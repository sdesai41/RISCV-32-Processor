
module datapath(clk);

input clk;
reg [11:0] PCnew,PCout,PCout2,PCim,PC4;
reg [11:0] PCresult,PCresultout;
reg [31:0]instruction,instrout;
reg signed [31:0] imm,immout;
reg [4:0] rs1,rs2,rd,rdout,rdo2,rdo3,rs1out,rs2out;
reg [31:0] op2;
reg signed [31:0] wdata;
reg signed [31:0] data1,data1out,data2,data2out,data2out2;
reg signed [31:0] op1fin,op2fin,data2fin;
reg pcsrc;
reg signed [31:0] result,resultout,resulto2,rdata, rdataout;
reg zero,neg;
reg zeroout,negout;
reg[4:0] aluop,aluopout,aluopu;
reg alusrc,alusrcout,alusrcu,memtoreg,memtoregu,memtoregout,memtorego2, memtorego3, regwrite,regwriteu,regwriteout,regwriteo2,regwriteo3,memreadu,memread,memwrite,memwriteu,sign,signu,signout,signout2,memwriteout,memwriteout2,memreadout,memreadout2;//sign for loads if we r signextending
reg [2:0] branch,branchout,branchout2,branchu;
reg [1:0] length,lengthout,lengthout2,lengthu;
reg ctrlf,pcwrite,fdwrite;
reg [1:0] forwardA,forwardB,forwardC;


initial begin 
PCim=0; 
pcsrc=0;
pcwrite=1;
fdwrite=1;
ctrlf=0;
forwardA=0;
forwardB=0;
forwardC=0;
end

add4 pcadd4(PCim,PC4);

instructionmemory IM(PCim,instruction);

fetchdecode reg1(clk,instruction, PCim,instrout,PCout, fdwrite);

decoder decode(instrout, rs1,rs2,rd,imm);

registerfile rf(rs1,rs2,rdo3,regwriteo3, wdata,data1,data2);

controller control(instrout, aluop,alusrc, memtoreg, regwrite,branch, memread,memwrite, length,sign );

controllermux flushctrl(ctrlf, aluop,alusrc, memtoreg, regwrite,branch,memread,memwrite,length,sign,aluopu,alusrcu, memtoregu, regwriteu,branchu,memreadu,memwriteu,lengthu,signu);

decodeex reg2(clk,rs1,rs1out,rs2,rs2out,PCout,imm,immout,data1,data2,rd,regwriteu,signu,memtoregu,memwriteu,memreadu,lengthu, alusrcu,branchu,aluopu,PCout2,data1out,data2out,rdout,regwriteout,signout,memtoregout,memreadout,lengthout, alusrcout,branchout,aluopout,memwriteout);

mux32 aluselect(immout,data2out,op2,alusrcout);

threemux32 aluforwardA(data1out,resultout,wdata,op1fin,forwardA);

threemux32 aluforwardB(op2,resultout,wdata,op2fin,forwardB); 

threemux32 data2forward(data2out, resultout,wdata,data2fin,forwardC);

ALU aluex(aluopout,signout,op1fin,op2fin,result,zero,neg);

pcadder PCADD(PCout2, immout, PCresult);

exmem reg3(clk,data2fin,data2out2,result,resultout,zero,zeroout,neg,negout,rdout,rdo2,PCresult, PCresultout, memreadout,memreadout2,memwriteout,memwriteout2, lengthout, lengthout2, signout, signout2, regwriteout,regwriteo2, memtoregout,memtorego2,branchout,branchout2);

datamemory mem(data2out2, resultout, memreadout2,memwriteout2,lengthout2,rdata,signout2);

branchdecision branchchoice(branchout2,zeroout,negout,pcsrc);

memwb reg4(clk,resultout,resulto2,rdata,rdataout,rdo3,rdo2,memtorego2, regwriteo2,memtorego3,regwriteo3);

mux32 writeback(rdataout, resulto2,wdata, memtorego3);

mux11 pcmux(PCresultout,PC4,PCnew,pcsrc);

forwardingunit FU(rs1out,rs2out,rdo2,rdo3,regwriteo2,regwriteo3,memreadout,memwriteout, forwardA,forwardB,forwardC);

hazard_detection HD(memreadout, rs1,rs2,rdout, ctrlf,pcwrite,fdwrite);

PCreg regpc(PCnew,clk,PCim,pcwrite);




endmodule







