module instructionmemory(PCn,data_out);
parameter PCSIZE=16;

reg [7:0] im [0:4095];
//input clk;
input reg [PCSIZE-1:0] PCn;
output reg [31:0] data_out;

initial begin // setting instruction memory
//PC=0;
//r-type
/*
im[0]=8'd19; 
im[1]= 8'd6; 
im[2]=8'd80; 
im[3]=8'd0;

im[4]=8'd147;
im[5]= 8'd102; 
im[6]=8'd176; 
im[7]=8'd0;

im[8]=8'd51; 
im[9]= 8'd135; 
im[10]=8'd198; 
im[11]=8'd0;
//data_in={8'd51, 8'd135,8'd198,8'd0};
im[12]=8'd179; 
im[13]= 8'd135;
 im[14]=8'd198;
 im[15]=8'd64;
im[16]=8'd19; 
im[17]= 8'd120; 
im[18]=8'd7; 
im[19]=8'd1;
im[20]=8'd179; 
im[20+1]= 8'd104;
im[20+2]=8'd216;
im[20+3]=8'd0;
im[24]=8'd51; 
im[24+1]= 8'd9; 
im[24+2]=8'd216; 
im[24+3]=8'd0;
*/
////lw/sw
/*
im[0]=8'd19; im[1]= 8'd6; im[2]=8'd80; im[3]=8'd0;

im[4]=8'd147; im[4+1]= 8'd102; im[4+2]=8'd176; im[4+3]=8'd0;

im[8]=8'd35; im[8+1]= 8'd34; im[8+2]=8'd192; im[8+3]=8'd0;

im[12]=8'd35; im[12+1]= 8'd36; im[12+2]=8'd208; im[12+3]=8'd0;

im[16]=8'd19; im[16+1]= 8'd118; im[16+2]=8'd6; im[16+3]=8'd0;

im[20]=8'd3; im[20+1]= 8'd38; im[20+2]=8'd70; im[20+3]=8'd0;

//copied line
im[24]=8'd3; im[24+1]= 8'd38; im[24+2]=8'd64; im[24+3]=8'd0;

im[28]=8'd51; im[28+1]= 8'd135; im[28+2]=8'd198; im[28+3]=8'd0;

im[32]=8'd179; im[32+1]= 8'd246; im[32+2]=8'd6; im[32+3]=8'd0;

im[36]=8'd179; im[36+1]= 8'd135; im[36+2]=8'd198; im[36+3]=8'd64;

im[40]=8'd131; im[40+1]= 8'd38; im[40+2]=8'd128; im[40+3]=8'd0;

im[44]=8'd51; im[44+1]= 8'd136; im[44+2]=8'd198; im[44+3]=8'd64;

im[48]=8'd179; im[48+1]= 8'd8; im[48+2]=8'd248; im[48+3]=8'd64;

im[52]=8'd131; im[52+1]= 8'd38; im[52+2]=8'd128; im[52+3]=8'd0;

*/


//branch

//im[0]=8'd19; im[1]= 8'd6; im[2]=8'd80; im[3]=8'd0;
//
//im[4]=8'd99; im[4+1]= 8'd4; im[4+2]=8'd6; im[4+3]=8'd6;
//
//im[8]=8'd35; im[8+1]= 8'd34; im[8+2]=8'd192; im[8+3]=8'd0;
//
//im[12]=8'd147; im[12+1]= 8'd6; im[12+2]=8'd112; im[12+3]=8'd0;
//
//im[16]=8'd99; im[16+1]= 8'd4; im[16+2]=8'd198; im[16+3]=8'd0;
//
//im[20]=8'd147; im[20+1]= 8'd102; im[20+2]=8'd240; im[20+3]=8'd0;
//
//im[24]=8'd3; im[24+1]= 8'd39; im[24+2]=8'd64; im[24+3]=8'd0;
//
//im[28]=8'd179; im[28+1]= 8'd135; im[28+2]=8'd230; im[28+3]=8'd64;
//
//im[32]=8'd35; im[32+1]= 8'd36; im[32+2]=8'd240; im[32+3]=8'd00;
//
//im[36]=8'd19; im[36+1]= 8'd8; im[36+2]=8'd0; im[36+3]=8'd0;
//
//im[40]=8'd51; im[40+1]= 8'd8; im[40+2]=8'd6; im[40+3]=8'd1;
//
//im[44]=8'd19; im[44+1]= 8'd6; im[44+2]=8'd246; im[44+3]=8'd255;
//
//im[48]=8'd99; im[48+1]= 8'd14; im[48+2]=8'd6; im[51]=8'd2;
//
//im[52]=8'd227 ; im[52+1]= 8'd10; im[54]=8'd198; im[55]=8'd254;
////*/
//AUTOMOTIVE BASIC LARGE
im[0]= 8'h13;
im[1]= 8'h01;
im[2]= 8'h01;
im[3]= 8'hFE;
im[4]= 8'h23;
im[5]= 8'h2E;
im[6]= 8'h11;
im[7]= 8'h00;
im[8]= 8'h23;
im[9]= 8'h2C;
im[10]= 8'h81;
im[11]= 8'h00;
im[12]= 8'h13;
im[13]= 8'h04;
im[14]= 8'h01;
im[15]= 8'h02;
im[16]= 8'h23;
im[17]= 8'h2A;
im[18]= 8'hA4;
im[19]= 8'hFE;
im[20]= 8'h23;
im[21]= 8'h28;
im[22]= 8'hB4;
im[23]= 8'hFE;
im[24]= 8'h23;
im[25]= 8'h26;
im[26]= 8'hA4;
im[27]= 8'hFE;
im[28]= 8'h23;
im[29]= 8'h24;
im[30]= 8'hA4;
im[31]= 8'hFE;
im[32]= 8'h23;
im[33]= 8'h22;
im[34]= 8'hA4;
im[35]= 8'hFE;
im[36]= 8'h23;
im[37]= 8'h20;
im[38]= 8'hA4;
im[39]= 8'hFE;
im[40]= 8'h6F;
im[41]= 8'h00;
im[42]= 8'h40;
im[43]= 8'h00;
im[44]= 8'h83;
im[45]= 8'h25;
im[46]= 8'h04;
im[47]= 8'hFE;
im[48]= 8'h13;
im[49]= 8'h05;
im[50]= 8'hF0;
im[51]= 8'h01;
im[52]= 8'h63;
im[53]= 8'h46;
im[54]= 8'hB5;
im[55]= 8'h08;
im[56]= 8'h6F;
im[57]= 8'h00;
im[58]= 8'h40;
im[59]= 8'h00;
im[60]= 8'h03;
im[61]= 8'h25;
im[62]= 8'h84;
im[63]= 8'hFE;
im[64]= 8'h13;
im[65]= 8'h15;
im[66]= 8'h25;
im[67]= 8'h00;
im[68]= 8'h83;
im[69]= 8'h25;
im[70]= 8'h44;
im[71]= 8'hFF;
im[72]= 8'h93;
im[73]= 8'hD5;
im[74]= 8'hE5;
im[75]= 8'h01;
im[76]= 8'h33;
im[77]= 8'h65;
im[78]= 8'hB5;
im[79]= 8'h00;
im[80]= 8'h23;
im[81]= 8'h24;
im[82]= 8'hA4;
im[83]= 8'hFE;
im[84]= 8'h03;
im[85]= 8'h25;
im[86]= 8'h44;
im[87]= 8'hFF;
im[88]= 8'h13;
im[89]= 8'h15;
im[90]= 8'h25;
im[91]= 8'h00;
im[92]= 8'h23;
im[93]= 8'h2A;
im[94]= 8'hA4;
im[95]= 8'hFE;
im[96]= 8'h03;
im[97]= 8'h25;
im[98]= 8'hC4;
im[99]= 8'hFE;
im[100]= 8'h13;
im[101]= 8'h15;
im[102]= 8'h15;
im[103]= 8'h00;
im[104]= 8'h23;
im[105]= 8'h26;
im[106]= 8'hA4;
im[107]= 8'hFE;
im[108]= 8'h03;
im[109]= 8'h25;
im[110]= 8'hC4;
im[111]= 8'hFE;
im[112]= 8'h13;
im[113]= 8'h15;
im[114]= 8'h15;
im[115]= 8'h00;
im[116]= 8'h13;
im[117]= 8'h65;
im[118]= 8'h15;
im[119]= 8'h00;
im[120]= 8'h23;
im[121]= 8'h22;
im[122]= 8'hA4;
im[123]= 8'hFE;
im[124]= 8'h03;
im[125]= 8'h25;
im[126]= 8'h84;
im[127]= 8'hFE;
im[128]= 8'h83;
im[129]= 8'h25;
im[130]= 8'h44;
im[131]= 8'hFE;
im[132]= 8'h63;
im[133]= 8'h64;
im[134]= 8'hB5;
im[135]= 8'h02;
im[136]= 8'h6F;
im[137]= 8'h00;
im[138]= 8'h40;
im[139]= 8'h00;
im[140]= 8'h83;
im[141]= 8'h25;
im[142]= 8'h44;
im[143]= 8'hFE;
im[144]= 8'h03;
im[145]= 8'h25;
im[146]= 8'h84;
im[147]= 8'hFE;
im[148]= 8'h33;
im[149]= 8'h05;
im[150]= 8'hB5;
im[151]= 8'h40;
im[152]= 8'h23;
im[153]= 8'h24;
im[154]= 8'hA4;
im[155]= 8'hFE;
im[156]= 8'h03;
im[157]= 8'h25;
im[158]= 8'hC4;
im[159]= 8'hFE;
im[160]= 8'h13;
im[161]= 8'h05;
im[162]= 8'h15;
im[163]= 8'h00;
im[164]= 8'h23;
im[165]= 8'h26;
im[166]= 8'hA4;
im[167]= 8'hFE;
im[168]= 8'h6F;
im[169]= 8'h00;
im[170]= 8'h40;
im[171]= 8'h00;
im[172]= 8'h6F;
im[173]= 8'h00;
im[174]= 8'h40;
im[175]= 8'h00;
im[176]= 8'h03;
im[177]= 8'h25;
im[178]= 8'h04;
im[179]= 8'hFE;
im[180]= 8'h13;
im[181]= 8'h05;
im[182]= 8'h15;
im[183]= 8'h00;
im[184]= 8'h23;
im[185]= 8'h20;
im[186]= 8'hA4;
im[187]= 8'hFE;
im[188]= 8'h6F;
im[189]= 8'hF0;
im[190]= 8'h1F;
im[191]= 8'hF7;
im[192]= 8'h83;
im[193]= 8'h25;
im[194]= 8'h04;
im[195]= 8'hFF;
im[196]= 8'h03;
im[197]= 8'h25;
im[198]= 8'hC4;
im[199]= 8'hFE;
im[200]= 8'h23;
im[201]= 8'hA0;
im[202]= 8'hA5;
im[203]= 8'h00;
im[204]= 8'h03;
im[205]= 8'h24;
im[206]= 8'h81;
im[207]= 8'h01;
im[208]= 8'h83;
im[209]= 8'h20;
im[210]= 8'hC1;
im[211]= 8'h01;
im[212]= 8'h13;
im[213]= 8'h01;
im[214]= 8'h01;
im[215]= 8'h02;
im[216]= 8'h13;
im[217]= 8'h01;
im[218]= 8'h01;
im[219]= 8'h81;
im[220]= 8'h23;
im[221]= 8'h26;
im[222]= 8'h11;
im[223]= 8'h7E;
im[224]= 8'h23;
im[225]= 8'h24;
im[226]= 8'h81;
im[227]= 8'h7E;
im[228]= 8'h13;
im[229]= 8'h04;
im[230]= 8'h01;
im[231]= 8'h7F;
im[232]= 8'h13;
im[233]= 8'h01;
im[234]= 8'h01;
im[235]= 8'hEE;
im[236]= 8'h23;
im[237]= 8'h26;
im[238]= 8'hA4;
im[239]= 8'hFC;
im[240]= 8'h23;
im[241]= 8'h24;
im[242]= 8'hB4;
im[243]= 8'hFC;
im[244]= 8'h13;
im[245]= 8'h05;
im[246]= 8'h04;
im[247]= 8'hF5;
im[248]= 8'h03;
im[249]= 8'h25;
im[250]= 8'h04;
im[251]= 8'hF5;
im[252]= 8'h83;
im[253]= 8'h25;
im[254]= 8'h44;
im[255]= 8'hF5;
im[256]= 8'h03;
im[257]= 8'h26;
im[258]= 8'h84;
im[259]= 8'hF5;
im[260]= 8'h83;
im[261]= 8'h26;
im[262]= 8'hC4;
im[263]= 8'hF5;
im[264]= 8'h23;
im[265]= 8'h2E;
im[266]= 8'hD4;
im[267]= 8'hFA;
im[268]= 8'h23;
im[269]= 8'h2C;
im[270]= 8'hC4;
im[271]= 8'hFA;
im[272]= 8'h23;
im[273]= 8'h2A;
im[274]= 8'hB4;
im[275]= 8'hFA;
im[276]= 8'h23;
im[277]= 8'h28;
im[278]= 8'hA4;
im[279]= 8'hFA;
im[280]= 8'h13;
im[281]= 8'h05;
im[282]= 8'h04;
im[283]= 8'hF4;
im[284]= 8'h03;
im[285]= 8'h25;
im[286]= 8'h04;
im[287]= 8'hF4;
im[288]= 8'h83;
im[289]= 8'h25;
im[290]= 8'h44;
im[291]= 8'hF4;
im[292]= 8'h03;
im[293]= 8'h26;
im[294]= 8'h84;
im[295]= 8'hF4;
im[296]= 8'h83;
im[297]= 8'h26;
im[298]= 8'hC4;
im[299]= 8'hF4;
im[300]= 8'h23;
im[301]= 8'h26;
im[302]= 8'hD4;
im[303]= 8'hFA;
im[304]= 8'h23;
im[305]= 8'h24;
im[306]= 8'hC4;
im[307]= 8'hFA;
im[308]= 8'h23;
im[309]= 8'h22;
im[310]= 8'hB4;
im[311]= 8'hFA;
im[312]= 8'h23;
im[313]= 8'h20;
im[314]= 8'hA4;
im[315]= 8'hFA;
im[316]= 8'h13;
im[317]= 8'h05;
im[318]= 8'h04;
im[319]= 8'hF3;
im[320]= 8'h03;
im[321]= 8'h25;
im[322]= 8'h04;
im[323]= 8'hF3;
im[324]= 8'h83;
im[325]= 8'h25;
im[326]= 8'h44;
im[327]= 8'hF3;
im[328]= 8'h03;
im[329]= 8'h26;
im[330]= 8'h84;
im[331]= 8'hF3;
im[332]= 8'h83;
im[333]= 8'h26;
im[334]= 8'hC4;
im[335]= 8'hF3;
im[336]= 8'h23;
im[337]= 8'h2E;
im[338]= 8'hD4;
im[339]= 8'hF8;
im[340]= 8'h23;
im[341]= 8'h2C;
im[342]= 8'hC4;
im[343]= 8'hF8;
im[344]= 8'h23;
im[345]= 8'h2A;
im[346]= 8'hB4;
im[347]= 8'hF8;
im[348]= 8'h23;
im[349]= 8'h28;
im[350]= 8'hA4;
im[351]= 8'hF8;
im[352]= 8'h03;
im[353]= 8'h25;
im[354]= 8'h04;
im[355]= 8'hFB;
im[356]= 8'h83;
im[357]= 8'h25;
im[358]= 8'h44;
im[359]= 8'hFB;
im[360]= 8'h03;
im[361]= 8'h26;
im[362]= 8'h84;
im[363]= 8'hFB;
im[364]= 8'h83;
im[365]= 8'h26;
im[366]= 8'hC4;
im[367]= 8'hFB;
im[368]= 8'h23;
im[369]= 8'h26;
im[370]= 8'hD4;
im[371]= 8'hF0;
im[372]= 8'h23;
im[373]= 8'h24;
im[374]= 8'hC4;
im[375]= 8'hF0;
im[376]= 8'h23;
im[377]= 8'h22;
im[378]= 8'hB4;
im[379]= 8'hF0;
im[380]= 8'h23;
im[381]= 8'h20;
im[382]= 8'hA4;
im[383]= 8'hF0;
im[384]= 8'h23;
im[385]= 8'h2E;
im[386]= 8'hD4;
im[387]= 8'hF0;
im[388]= 8'h23;
im[389]= 8'h2C;
im[390]= 8'hC4;
im[391]= 8'hF0;
im[392]= 8'h23;
im[393]= 8'h2A;
im[394]= 8'hB4;
im[395]= 8'hF0;
im[396]= 8'h23;
im[397]= 8'h28;
im[398]= 8'hA4;
im[399]= 8'hF0;
im[400]= 8'h13;
im[401]= 8'h05;
im[402]= 8'h04;
im[403]= 8'hF2;
im[404]= 8'h93;
im[405]= 8'h05;
im[406]= 8'h04;
im[407]= 8'hF1;
im[408]= 8'h13;
im[409]= 8'h06;
im[410]= 8'h04;
im[411]= 8'hF0;
im[412]= 8'h03;
im[413]= 8'h25;
im[414]= 8'h04;
im[415]= 8'hF2;
im[416]= 8'h93;
im[417]= 8'h85;
im[418]= 8'h45;
im[419]= 8'h7F;
im[420]= 8'hB3;
im[421]= 8'h85;
im[422]= 8'h85;
im[423]= 8'h00;
im[424]= 8'h23;
im[425]= 8'hA0;
im[426]= 8'hA5;
im[427]= 8'h00;
im[428]= 8'h03;
im[429]= 8'h25;
im[430]= 8'h44;
im[431]= 8'hF2;
im[432]= 8'h93;
im[433]= 8'h85;
im[434]= 8'h05;
im[435]= 8'h7F;
im[436]= 8'hB3;
im[437]= 8'h85;
im[438]= 8'h85;
im[439]= 8'h00;
im[440]= 8'h23;
im[441]= 8'hA0;
im[442]= 8'hA5;
im[443]= 8'h00;
im[444]= 8'h03;
im[445]= 8'h25;
im[446]= 8'h84;
im[447]= 8'hF2;
im[448]= 8'h93;
im[449]= 8'h85;
im[450]= 8'hC5;
im[451]= 8'h7E;
im[452]= 8'hB3;
im[453]= 8'h85;
im[454]= 8'h85;
im[455]= 8'h00;
im[456]= 8'h23;
im[457]= 8'hA0;
im[458]= 8'hA5;
im[459]= 8'h00;
im[460]= 8'h03;
im[461]= 8'h25;
im[462]= 8'hC4;
im[463]= 8'hF2;
im[464]= 8'h93;
im[465]= 8'h85;
im[466]= 8'h85;
im[467]= 8'h7E;
im[468]= 8'hB3;
im[469]= 8'h85;
im[470]= 8'h85;
im[471]= 8'h00;
im[472]= 8'h23;
im[473]= 8'hA0;
im[474]= 8'hA5;
im[475]= 8'h00;
im[476]= 8'h03;
im[477]= 8'h25;
im[478]= 8'h04;
im[479]= 8'hFA;
im[480]= 8'h83;
im[481]= 8'h25;
im[482]= 8'h44;
im[483]= 8'hFA;
im[484]= 8'h03;
im[485]= 8'h26;
im[486]= 8'h84;
im[487]= 8'hFA;
im[488]= 8'h83;
im[489]= 8'h26;
im[490]= 8'hC4;
im[491]= 8'hFA;
im[492]= 8'h23;
im[493]= 8'h2E;
im[494]= 8'hE4;
im[495]= 8'hEC;
im[496]= 8'h23;
im[497]= 8'h26;
im[498]= 8'hE4;
im[499]= 8'h82;
im[500]= 8'h23;
im[501]= 8'h2C;
im[502]= 8'hE4;
im[503]= 8'hEC;
im[504]= 8'h23;
im[505]= 8'h2A;
im[506]= 8'hE4;
im[507]= 8'hEC;
im[508]= 8'h23;
im[509]= 8'h28;
im[510]= 8'hE4;
im[511]= 8'hEC;
im[512]= 8'h23;
im[513]= 8'h26;
im[514]= 8'hD4;
im[515]= 8'hEE;
im[516]= 8'h23;
im[517]= 8'h24;
im[518]= 8'hC4;
im[519]= 8'hEE;
im[520]= 8'h23;
im[521]= 8'h22;
im[522]= 8'hB4;
im[523]= 8'hEE;
im[524]= 8'h23;
im[525]= 8'h20;
im[526]= 8'hA4;
im[527]= 8'hEE;
im[528]= 8'h13;
im[529]= 8'h05;
im[530]= 8'h04;
im[531]= 8'hEF;
im[532]= 8'h93;
im[533]= 8'h05;
im[534]= 8'h04;
im[535]= 8'hEE;
im[536]= 8'h13;
im[537]= 8'h06;
im[538]= 8'h04;
im[539]= 8'hED;
im[540]= 8'h13;
im[541]= 8'h05;
im[542]= 8'h85;
im[543]= 8'h7E;
im[544]= 8'h33;
im[545]= 8'h05;
im[546]= 8'h85;
im[547]= 8'h00;
im[548]= 8'h83;
im[549]= 8'h26;
im[550]= 8'h05;
im[551]= 8'h00;
im[552]= 8'h13;
im[553]= 8'h05;
im[554]= 8'hC5;
im[555]= 8'h7E;
im[556]= 8'h33;
im[557]= 8'h05;
im[558]= 8'h85;
im[559]= 8'h00;
im[560]= 8'h03;
im[561]= 8'h26;
im[562]= 8'h05;
im[563]= 8'h00;
im[564]= 8'h13;
im[565]= 8'h05;
im[566]= 8'h05;
im[567]= 8'h7F;
im[568]= 8'h33;
im[569]= 8'h05;
im[570]= 8'h85;
im[571]= 8'h00;
im[572]= 8'h83;
im[573]= 8'h25;
im[574]= 8'h05;
im[575]= 8'h00;
im[576]= 8'h13;
im[577]= 8'h05;
im[578]= 8'h45;
im[579]= 8'h7F;
im[580]= 8'h33;
im[581]= 8'h05;
im[582]= 8'h85;
im[583]= 8'h00;
im[584]= 8'h03;
im[585]= 8'h25;
im[586]= 8'h05;
im[587]= 8'h00;
im[588]= 8'h03;
im[589]= 8'h27;
im[590]= 8'h04;
im[591]= 8'hEF;
im[592]= 8'h83;
im[593]= 8'h27;
im[594]= 8'h44;
im[595]= 8'hEF;
im[596]= 8'h03;
im[597]= 8'h28;
im[598]= 8'h84;
im[599]= 8'hEF;
im[600]= 8'h83;
im[601]= 8'h28;
im[602]= 8'hC4;
im[603]= 8'hEF;
im[604]= 8'h23;
im[605]= 8'h26;
im[606]= 8'h14;
im[607]= 8'hEB;
im[608]= 8'h23;
im[609]= 8'h24;
im[610]= 8'h04;
im[611]= 8'hEB;
im[612]= 8'h23;
im[613]= 8'h22;
im[614]= 8'hF4;
im[615]= 8'hEA;
im[616]= 8'h23;
im[617]= 8'h20;
im[618]= 8'hE4;
im[619]= 8'hEA;
im[620]= 8'h23;
im[621]= 8'h2E;
im[622]= 8'hD4;
im[623]= 8'hEA;
im[624]= 8'h23;
im[625]= 8'h2C;
im[626]= 8'hC4;
im[627]= 8'hEA;
im[628]= 8'h23;
im[629]= 8'h2A;
im[630]= 8'hB4;
im[631]= 8'hEA;
im[632]= 8'h23;
im[633]= 8'h28;
im[634]= 8'hA4;
im[635]= 8'hEA;
im[636]= 8'h13;
im[637]= 8'h05;
im[638]= 8'h04;
im[639]= 8'hEC;
im[640]= 8'h93;
im[641]= 8'h05;
im[642]= 8'h04;
im[643]= 8'hEB;
im[644]= 8'h13;
im[645]= 8'h06;
im[646]= 8'h04;
im[647]= 8'hEA;
im[648]= 8'h03;
im[649]= 8'h27;
im[650]= 8'hC4;
im[651]= 8'h82;
im[652]= 8'h03;
im[653]= 8'h25;
im[654]= 8'h04;
im[655]= 8'hEC;
im[656]= 8'h83;
im[657]= 8'h25;
im[658]= 8'h44;
im[659]= 8'hEC;
im[660]= 8'h03;
im[661]= 8'h26;
im[662]= 8'h84;
im[663]= 8'hEC;
im[664]= 8'h83;
im[665]= 8'h26;
im[666]= 8'hC4;
im[667]= 8'hEC;
im[668]= 8'h13;
im[669]= 8'h08;
im[670]= 8'h88;
im[671]= 8'h7F;
im[672]= 8'h33;
im[673]= 8'h08;
im[674]= 8'h88;
im[675]= 8'h00;
im[676]= 8'h23;
im[677]= 8'h20;
im[678]= 8'hF8;
im[679]= 8'h00;
im[680]= 8'h23;
im[681]= 8'h2E;
im[682]= 8'hF4;
im[683]= 8'hE6;
im[684]= 8'h23;
im[685]= 8'h2C;
im[686]= 8'hE4;
im[687]= 8'hE6;
im[688]= 8'h23;
im[689]= 8'h2A;
im[690]= 8'hE4;
im[691]= 8'hE6;
im[692]= 8'h23;
im[693]= 8'h28;
im[694]= 8'hE4;
im[695]= 8'hE6;
im[696]= 8'h23;
im[697]= 8'h26;
im[698]= 8'hD4;
im[699]= 8'hE8;
im[700]= 8'h23;
im[701]= 8'h24;
im[702]= 8'hC4;
im[703]= 8'hE8;
im[704]= 8'h23;
im[705]= 8'h22;
im[706]= 8'hB4;
im[707]= 8'hE8;
im[708]= 8'h23;
im[709]= 8'h20;
im[710]= 8'hA4;
im[711]= 8'hE8;
im[712]= 8'h13;
im[713]= 8'h05;
im[714]= 8'h04;
im[715]= 8'hE9;
im[716]= 8'h93;
im[717]= 8'h05;
im[718]= 8'h04;
im[719]= 8'hE8;
im[720]= 8'h13;
im[721]= 8'h06;
im[722]= 8'h04;
im[723]= 8'hE7;
im[724]= 8'h03;
im[725]= 8'h25;
im[726]= 8'h04;
im[727]= 8'hE9;
im[728]= 8'h83;
im[729]= 8'h25;
im[730]= 8'h44;
im[731]= 8'hE9;
im[732]= 8'h03;
im[733]= 8'h26;
im[734]= 8'h84;
im[735]= 8'hE9;
im[736]= 8'h83;
im[737]= 8'h26;
im[738]= 8'hC4;
im[739]= 8'hE9;
im[740]= 8'h23;
im[741]= 8'h26;
im[742]= 8'hD4;
im[743]= 8'hF8;
im[744]= 8'h23;
im[745]= 8'h24;
im[746]= 8'hC4;
im[747]= 8'hF8;
im[748]= 8'h23;
im[749]= 8'h22;
im[750]= 8'hB4;
im[751]= 8'hF8;
im[752]= 8'h23;
im[753]= 8'h20;
im[754]= 8'hA4;
im[755]= 8'hF8;
im[756]= 8'h03;
im[757]= 8'h25;
im[758]= 8'h04;
im[759]= 8'hFB;
im[760]= 8'h23;
im[761]= 8'h24;
im[762]= 8'hA4;
im[763]= 8'h80;
im[764]= 8'h83;
im[765]= 8'h25;
im[766]= 8'h44;
im[767]= 8'hFB;
im[768]= 8'h23;
im[769]= 8'h22;
im[770]= 8'hB4;
im[771]= 8'h80;
im[772]= 8'h03;
im[773]= 8'h26;
im[774]= 8'h84;
im[775]= 8'hFB;
im[776]= 8'h23;
im[777]= 8'h20;
im[778]= 8'hC4;
im[779]= 8'h80;
im[780]= 8'h83;
im[781]= 8'h26;
im[782]= 8'hC4;
im[783]= 8'hFB;
im[784]= 8'h13;
im[785]= 8'h07;
im[786]= 8'hC7;
im[787]= 8'h7F;
im[788]= 8'h33;
im[789]= 8'h07;
im[790]= 8'h87;
im[791]= 8'h00;
im[792]= 8'h23;
im[793]= 8'h20;
im[794]= 8'hD7;
im[795]= 8'h00;
im[796]= 8'h23;
im[797]= 8'h2E;
im[798]= 8'hD4;
im[799]= 8'hE0;
im[800]= 8'h23;
im[801]= 8'h2C;
im[802]= 8'hC4;
im[803]= 8'hE0;
im[804]= 8'h23;
im[805]= 8'h2A;
im[806]= 8'hB4;
im[807]= 8'hE0;
im[808]= 8'h23;
im[809]= 8'h28;
im[810]= 8'hA4;
im[811]= 8'hE0;
im[812]= 8'h23;
im[813]= 8'h26;
im[814]= 8'hD4;
im[815]= 8'hE2;
im[816]= 8'h23;
im[817]= 8'h24;
im[818]= 8'hC4;
im[819]= 8'hE2;
im[820]= 8'h23;
im[821]= 8'h22;
im[822]= 8'hB4;
im[823]= 8'hE2;
im[824]= 8'h23;
im[825]= 8'h20;
im[826]= 8'hA4;
im[827]= 8'hE2;
im[828]= 8'h13;
im[829]= 8'h05;
im[830]= 8'h04;
im[831]= 8'hE3;
im[832]= 8'h93;
im[833]= 8'h05;
im[834]= 8'h04;
im[835]= 8'hE2;
im[836]= 8'h13;
im[837]= 8'h06;
im[838]= 8'h04;
im[839]= 8'hE1;
im[840]= 8'h13;
im[841]= 8'h05;
im[842]= 8'hC5;
im[843]= 8'h7F;
im[844]= 8'h33;
im[845]= 8'h05;
im[846]= 8'h85;
im[847]= 8'h00;
im[848]= 8'h83;
im[849]= 8'h28;
im[850]= 8'h05;
im[851]= 8'h00;
im[852]= 8'h03;
im[853]= 8'h28;
im[854]= 8'h04;
im[855]= 8'h80;
im[856]= 8'h83;
im[857]= 8'h27;
im[858]= 8'h44;
im[859]= 8'h80;
im[860]= 8'h03;
im[861]= 8'h27;
im[862]= 8'h84;
im[863]= 8'h80;
im[864]= 8'h03;
im[865]= 8'h25;
im[866]= 8'h04;
im[867]= 8'hE3;
im[868]= 8'h83;
im[869]= 8'h25;
im[870]= 8'h44;
im[871]= 8'hE3;
im[872]= 8'h03;
im[873]= 8'h26;
im[874]= 8'h84;
im[875]= 8'hE3;
im[876]= 8'h83;
im[877]= 8'h26;
im[878]= 8'hC4;
im[879]= 8'hE3;
im[880]= 8'h23;
im[881]= 8'h26;
im[882]= 8'h14;
im[883]= 8'hDF;
im[884]= 8'h23;
im[885]= 8'h24;
im[886]= 8'h04;
im[887]= 8'hDF;
im[888]= 8'h23;
im[889]= 8'h22;
im[890]= 8'hF4;
im[891]= 8'hDE;
im[892]= 8'h23;
im[893]= 8'h20;
im[894]= 8'hE4;
im[895]= 8'hDE;
im[896]= 8'h23;
im[897]= 8'h2E;
im[898]= 8'hD4;
im[899]= 8'hDE;
im[900]= 8'h23;
im[901]= 8'h2C;
im[902]= 8'hC4;
im[903]= 8'hDE;
im[904]= 8'h23;
im[905]= 8'h2A;
im[906]= 8'hB4;
im[907]= 8'hDE;
im[908]= 8'h23;
im[909]= 8'h28;
im[910]= 8'hA4;
im[911]= 8'hDE;
im[912]= 8'h13;
im[913]= 8'h05;
im[914]= 8'h04;
im[915]= 8'hE0;
im[916]= 8'h93;
im[917]= 8'h05;
im[918]= 8'h04;
im[919]= 8'hDF;
im[920]= 8'h13;
im[921]= 8'h06;
im[922]= 8'h04;
im[923]= 8'hDE;
im[924]= 8'h13;
im[925]= 8'h05;
im[926]= 8'hC5;
im[927]= 8'h7F;
im[928]= 8'h33;
im[929]= 8'h05;
im[930]= 8'h85;
im[931]= 8'h00;
im[932]= 8'h83;
im[933]= 8'h28;
im[934]= 8'h05;
im[935]= 8'h00;
im[936]= 8'h03;
im[937]= 8'h28;
im[938]= 8'h04;
im[939]= 8'h80;
im[940]= 8'h83;
im[941]= 8'h27;
im[942]= 8'h44;
im[943]= 8'h80;
im[944]= 8'h03;
im[945]= 8'h27;
im[946]= 8'h84;
im[947]= 8'h80;
im[948]= 8'h03;
im[949]= 8'h25;
im[950]= 8'h04;
im[951]= 8'hE0;
im[952]= 8'h83;
im[953]= 8'h25;
im[954]= 8'h44;
im[955]= 8'hE0;
im[956]= 8'h03;
im[957]= 8'h26;
im[958]= 8'h84;
im[959]= 8'hE0;
im[960]= 8'h83;
im[961]= 8'h26;
im[962]= 8'hC4;
im[963]= 8'hE0;
im[964]= 8'h23;
im[965]= 8'h2E;
im[966]= 8'h14;
im[967]= 8'hDB;
im[968]= 8'h23;
im[969]= 8'h2C;
im[970]= 8'h04;
im[971]= 8'hDB;
im[972]= 8'h23;
im[973]= 8'h2A;
im[974]= 8'hF4;
im[975]= 8'hDA;
im[976]= 8'h23;
im[977]= 8'h28;
im[978]= 8'hE4;
im[979]= 8'hDA;
im[980]= 8'h23;
im[981]= 8'h26;
im[982]= 8'hD4;
im[983]= 8'hDC;
im[984]= 8'h23;
im[985]= 8'h24;
im[986]= 8'hC4;
im[987]= 8'hDC;
im[988]= 8'h23;
im[989]= 8'h22;
im[990]= 8'hB4;
im[991]= 8'hDC;
im[992]= 8'h23;
im[993]= 8'h20;
im[994]= 8'hA4;
im[995]= 8'hDC;
im[996]= 8'h13;
im[997]= 8'h05;
im[998]= 8'h04;
im[999]= 8'hDD;
im[1000]= 8'h93;
im[1001]= 8'h05;
im[1002]= 8'h04;
im[1003]= 8'hDC;
im[1004]= 8'h13;
im[1005]= 8'h06;
im[1006]= 8'h04;
im[1007]= 8'hDB;
im[1008]= 8'h13;
im[1009]= 8'h05;
im[1010]= 8'h85;
im[1011]= 8'h7F;
im[1012]= 8'h33;
im[1013]= 8'h05;
im[1014]= 8'h85;
im[1015]= 8'h00;
im[1016]= 8'h83;
im[1017]= 8'h27;
im[1018]= 8'h05;
im[1019]= 8'h00;
im[1020]= 8'h13;
im[1021]= 8'h05;
im[1022]= 8'hC5;
im[1023]= 8'h7F;
im[1024]= 8'h33;
im[1025]= 8'h05;
im[1026]= 8'h85;
im[1027]= 8'h00;
im[1028]= 8'h83;
im[1029]= 8'h26;
im[1030]= 8'h05;
im[1031]= 8'h00;
im[1032]= 8'h03;
im[1033]= 8'h26;
im[1034]= 8'h04;
im[1035]= 8'h80;
im[1036]= 8'h83;
im[1037]= 8'h25;
im[1038]= 8'h44;
im[1039]= 8'h80;
im[1040]= 8'h03;
im[1041]= 8'h25;
im[1042]= 8'h84;
im[1043]= 8'h80;
im[1044]= 8'h03;
im[1045]= 8'h27;
im[1046]= 8'hC4;
im[1047]= 8'h82;
im[1048]= 8'h03;
im[1049]= 8'h28;
im[1050]= 8'h04;
im[1051]= 8'hDD;
im[1052]= 8'h23;
im[1053]= 8'h2C;
im[1054]= 8'h04;
im[1055]= 8'h81;
im[1056]= 8'h03;
im[1057]= 8'h28;
im[1058]= 8'h44;
im[1059]= 8'hDD;
im[1060]= 8'h23;
im[1061]= 8'h2A;
im[1062]= 8'h04;
im[1063]= 8'h81;
im[1064]= 8'h03;
im[1065]= 8'h28;
im[1066]= 8'h84;
im[1067]= 8'hDD;
im[1068]= 8'h23;
im[1069]= 8'h28;
im[1070]= 8'h04;
im[1071]= 8'h81;
im[1072]= 8'h03;
im[1073]= 8'h28;
im[1074]= 8'hC4;
im[1075]= 8'hDD;
im[1076]= 8'h23;
im[1077]= 8'h26;
im[1078]= 8'h04;
im[1079]= 8'h81;
im[1080]= 8'h23;
im[1081]= 8'h26;
im[1082]= 8'hF4;
im[1083]= 8'hE4;
im[1084]= 8'h23;
im[1085]= 8'h24;
im[1086]= 8'hE4;
im[1087]= 8'hE4;
im[1088]= 8'h23;
im[1089]= 8'h22;
im[1090]= 8'hE4;
im[1091]= 8'hE4;
im[1092]= 8'h23;
im[1093]= 8'h20;
im[1094]= 8'hE4;
im[1095]= 8'hE4;
im[1096]= 8'h23;
im[1097]= 8'h2E;
im[1098]= 8'hD4;
im[1099]= 8'hE4;
im[1100]= 8'h23;
im[1101]= 8'h2C;
im[1102]= 8'hC4;
im[1103]= 8'hE4;
im[1104]= 8'h23;
im[1105]= 8'h2A;
im[1106]= 8'hB4;
im[1107]= 8'hE4;
im[1108]= 8'h23;
im[1109]= 8'h28;
im[1110]= 8'hA4;
im[1111]= 8'hE4;
im[1112]= 8'h13;
im[1113]= 8'h05;
im[1114]= 8'h04;
im[1115]= 8'hE6;
im[1116]= 8'h93;
im[1117]= 8'h05;
im[1118]= 8'h04;
im[1119]= 8'hE5;
im[1120]= 8'h13;
im[1121]= 8'h06;
im[1122]= 8'h04;
im[1123]= 8'hE4;
im[1124]= 8'h03;
im[1125]= 8'h25;
im[1126]= 8'h04;
im[1127]= 8'hE6;
im[1128]= 8'h83;
im[1129]= 8'h25;
im[1130]= 8'h44;
im[1131]= 8'hE6;
im[1132]= 8'h03;
im[1133]= 8'h26;
im[1134]= 8'h84;
im[1135]= 8'hE6;
im[1136]= 8'h83;
im[1137]= 8'h26;
im[1138]= 8'hC4;
im[1139]= 8'hE6;
im[1140]= 8'h03;
im[1141]= 8'h27;
im[1142]= 8'h04;
im[1143]= 8'hFA;
im[1144]= 8'h83;
im[1145]= 8'h27;
im[1146]= 8'h44;
im[1147]= 8'hFA;
im[1148]= 8'h03;
im[1149]= 8'h28;
im[1150]= 8'h84;
im[1151]= 8'hFA;
im[1152]= 8'h83;
im[1153]= 8'h28;
im[1154]= 8'hC4;
im[1155]= 8'hFA;
im[1156]= 8'h23;
im[1157]= 8'h26;
im[1158]= 8'h14;
im[1159]= 8'hD9;
im[1160]= 8'h23;
im[1161]= 8'h24;
im[1162]= 8'h04;
im[1163]= 8'hD9;
im[1164]= 8'h23;
im[1165]= 8'h22;
im[1166]= 8'hF4;
im[1167]= 8'hD8;
im[1168]= 8'h23;
im[1169]= 8'h20;
im[1170]= 8'hE4;
im[1171]= 8'hD8;
im[1172]= 8'h23;
im[1173]= 8'h2E;
im[1174]= 8'hD4;
im[1175]= 8'hD8;
im[1176]= 8'h23;
im[1177]= 8'h2C;
im[1178]= 8'hC4;
im[1179]= 8'hD8;
im[1180]= 8'h23;
im[1181]= 8'h2A;
im[1182]= 8'hB4;
im[1183]= 8'hD8;
im[1184]= 8'h23;
im[1185]= 8'h28;
im[1186]= 8'hA4;
im[1187]= 8'hD8;
im[1188]= 8'h13;
im[1189]= 8'h05;
im[1190]= 8'h04;
im[1191]= 8'hDA;
im[1192]= 8'h93;
im[1193]= 8'h05;
im[1194]= 8'h04;
im[1195]= 8'hD9;
im[1196]= 8'h13;
im[1197]= 8'h06;
im[1198]= 8'h04;
im[1199]= 8'hD8;
im[1200]= 8'h83;
im[1201]= 8'h26;
im[1202]= 8'hC4;
im[1203]= 8'h80;
im[1204]= 8'h03;
im[1205]= 8'h26;
im[1206]= 8'h04;
im[1207]= 8'h81;
im[1208]= 8'h83;
im[1209]= 8'h25;
im[1210]= 8'h44;
im[1211]= 8'h81;
im[1212]= 8'h03;
im[1213]= 8'h25;
im[1214]= 8'h84;
im[1215]= 8'h81;
im[1216]= 8'h03;
im[1217]= 8'h27;
im[1218]= 8'h04;
im[1219]= 8'hDA;
im[1220]= 8'h83;
im[1221]= 8'h27;
im[1222]= 8'h44;
im[1223]= 8'hDA;
im[1224]= 8'h03;
im[1225]= 8'h28;
im[1226]= 8'h84;
im[1227]= 8'hDA;
im[1228]= 8'h83;
im[1229]= 8'h28;
im[1230]= 8'hC4;
im[1231]= 8'hDA;
im[1232]= 8'h23;
im[1233]= 8'h2E;
im[1234]= 8'h14;
im[1235]= 8'hD5;
im[1236]= 8'h23;
im[1237]= 8'h2C;
im[1238]= 8'h04;
im[1239]= 8'hD5;
im[1240]= 8'h23;
im[1241]= 8'h2A;
im[1242]= 8'hF4;
im[1243]= 8'hD4;
im[1244]= 8'h23;
im[1245]= 8'h28;
im[1246]= 8'hE4;
im[1247]= 8'hD4;
im[1248]= 8'h23;
im[1249]= 8'h26;
im[1250]= 8'hD4;
im[1251]= 8'hD6;
im[1252]= 8'h23;
im[1253]= 8'h24;
im[1254]= 8'hC4;
im[1255]= 8'hD6;
im[1256]= 8'h23;
im[1257]= 8'h22;
im[1258]= 8'hB4;
im[1259]= 8'hD6;
im[1260]= 8'h23;
im[1261]= 8'h20;
im[1262]= 8'hA4;
im[1263]= 8'hD6;
im[1264]= 8'h13;
im[1265]= 8'h05;
im[1266]= 8'h04;
im[1267]= 8'hD7;
im[1268]= 8'h93;
im[1269]= 8'h05;
im[1270]= 8'h04;
im[1271]= 8'hD6;
im[1272]= 8'h13;
im[1273]= 8'h06;
im[1274]= 8'h04;
im[1275]= 8'hD5;
im[1276]= 8'h03;
im[1277]= 8'h27;
im[1278]= 8'hC4;
im[1279]= 8'h82;
im[1280]= 8'h03;
im[1281]= 8'h25;
im[1282]= 8'h04;
im[1283]= 8'hD7;
im[1284]= 8'h23;
im[1285]= 8'h24;
im[1286]= 8'hA4;
im[1287]= 8'h82;
im[1288]= 8'h03;
im[1289]= 8'h25;
im[1290]= 8'h44;
im[1291]= 8'hD7;
im[1292]= 8'h23;
im[1293]= 8'h22;
im[1294]= 8'hA4;
im[1295]= 8'h82;
im[1296]= 8'h03;
im[1297]= 8'h25;
im[1298]= 8'h84;
im[1299]= 8'hD7;
im[1300]= 8'h23;
im[1301]= 8'h20;
im[1302]= 8'hA4;
im[1303]= 8'h82;
im[1304]= 8'h03;
im[1305]= 8'h25;
im[1306]= 8'hC4;
im[1307]= 8'hD7;
im[1308]= 8'h23;
im[1309]= 8'h2E;
im[1310]= 8'hA4;
im[1311]= 8'h80;
im[1312]= 8'h03;
im[1313]= 8'h25;
im[1314]= 8'h04;
im[1315]= 8'hF9;
im[1316]= 8'h83;
im[1317]= 8'h25;
im[1318]= 8'h44;
im[1319]= 8'hF9;
im[1320]= 8'h03;
im[1321]= 8'h26;
im[1322]= 8'h84;
im[1323]= 8'hF9;
im[1324]= 8'h83;
im[1325]= 8'h26;
im[1326]= 8'hC4;
im[1327]= 8'hF9;
im[1328]= 8'h23;
im[1329]= 8'h26;
im[1330]= 8'hF4;
im[1331]= 8'hD2;
im[1332]= 8'h23;
im[1333]= 8'h24;
im[1334]= 8'hE4;
im[1335]= 8'hD2;
im[1336]= 8'h23;
im[1337]= 8'h22;
im[1338]= 8'hE4;
im[1339]= 8'hD2;
im[1340]= 8'h23;
im[1341]= 8'h20;
im[1342]= 8'hE4;
im[1343]= 8'hD2;
im[1344]= 8'h23;
im[1345]= 8'h2E;
im[1346]= 8'hD4;
im[1347]= 8'hD2;
im[1348]= 8'h23;
im[1349]= 8'h2C;
im[1350]= 8'hC4;
im[1351]= 8'hD2;
im[1352]= 8'h23;
im[1353]= 8'h2A;
im[1354]= 8'hB4;
im[1355]= 8'hD2;
im[1356]= 8'h23;
im[1357]= 8'h28;
im[1358]= 8'hA4;
im[1359]= 8'hD2;
im[1360]= 8'h13;
im[1361]= 8'h05;
im[1362]= 8'h04;
im[1363]= 8'hD4;
im[1364]= 8'h93;
im[1365]= 8'h05;
im[1366]= 8'h04;
im[1367]= 8'hD3;
im[1368]= 8'h13;
im[1369]= 8'h06;
im[1370]= 8'h04;
im[1371]= 8'hD2;
im[1372]= 8'h83;
im[1373]= 8'h26;
im[1374]= 8'hC4;
im[1375]= 8'h81;
im[1376]= 8'h03;
im[1377]= 8'h26;
im[1378]= 8'h04;
im[1379]= 8'h82;
im[1380]= 8'h83;
im[1381]= 8'h25;
im[1382]= 8'h44;
im[1383]= 8'h82;
im[1384]= 8'h03;
im[1385]= 8'h25;
im[1386]= 8'h84;
im[1387]= 8'h82;
im[1388]= 8'h03;
im[1389]= 8'h27;
im[1390]= 8'h04;
im[1391]= 8'hD4;
im[1392]= 8'h83;
im[1393]= 8'h27;
im[1394]= 8'h44;
im[1395]= 8'hD4;
im[1396]= 8'h03;
im[1397]= 8'h28;
im[1398]= 8'h84;
im[1399]= 8'hD4;
im[1400]= 8'h83;
im[1401]= 8'h28;
im[1402]= 8'hC4;
im[1403]= 8'hD4;
im[1404]= 8'h23;
im[1405]= 8'h2E;
im[1406]= 8'h14;
im[1407]= 8'hCF;
im[1408]= 8'h23;
im[1409]= 8'h2C;
im[1410]= 8'h04;
im[1411]= 8'hCF;
im[1412]= 8'h23;
im[1413]= 8'h2A;
im[1414]= 8'hF4;
im[1415]= 8'hCE;
im[1416]= 8'h23;
im[1417]= 8'h28;
im[1418]= 8'hE4;
im[1419]= 8'hCE;
im[1420]= 8'h23;
im[1421]= 8'h26;
im[1422]= 8'hD4;
im[1423]= 8'hD0;
im[1424]= 8'h23;
im[1425]= 8'h24;
im[1426]= 8'hC4;
im[1427]= 8'hD0;
im[1428]= 8'h23;
im[1429]= 8'h22;
im[1430]= 8'hB4;
im[1431]= 8'hD0;
im[1432]= 8'h23;
im[1433]= 8'h20;
im[1434]= 8'hA4;
im[1435]= 8'hD0;
im[1436]= 8'h13;
im[1437]= 8'h05;
im[1438]= 8'h04;
im[1439]= 8'hD1;
im[1440]= 8'h93;
im[1441]= 8'h05;
im[1442]= 8'h04;
im[1443]= 8'hD0;
im[1444]= 8'h13;
im[1445]= 8'h06;
im[1446]= 8'h04;
im[1447]= 8'hCF;
im[1448]= 8'h03;
im[1449]= 8'h27;
im[1450]= 8'hC4;
im[1451]= 8'h82;
im[1452]= 8'h03;
im[1453]= 8'h25;
im[1454]= 8'h04;
im[1455]= 8'hD1;
im[1456]= 8'h83;
im[1457]= 8'h25;
im[1458]= 8'h44;
im[1459]= 8'hD1;
im[1460]= 8'h03;
im[1461]= 8'h26;
im[1462]= 8'h84;
im[1463]= 8'hD1;
im[1464]= 8'h83;
im[1465]= 8'h26;
im[1466]= 8'hC4;
im[1467]= 8'hD1;
im[1468]= 8'h23;
im[1469]= 8'h26;
im[1470]= 8'hF4;
im[1471]= 8'hCC;
im[1472]= 8'h23;
im[1473]= 8'h24;
im[1474]= 8'hE4;
im[1475]= 8'hCC;
im[1476]= 8'h23;
im[1477]= 8'h22;
im[1478]= 8'hE4;
im[1479]= 8'hCC;
im[1480]= 8'h23;
im[1481]= 8'h20;
im[1482]= 8'hE4;
im[1483]= 8'hCC;
im[1484]= 8'h23;
im[1485]= 8'h2E;
im[1486]= 8'hD4;
im[1487]= 8'hCC;
im[1488]= 8'h23;
im[1489]= 8'h2C;
im[1490]= 8'hC4;
im[1491]= 8'hCC;
im[1492]= 8'h23;
im[1493]= 8'h2A;
im[1494]= 8'hB4;
im[1495]= 8'hCC;
im[1496]= 8'h23;
im[1497]= 8'h28;
im[1498]= 8'hA4;
im[1499]= 8'hCC;
im[1500]= 8'h13;
im[1501]= 8'h05;
im[1502]= 8'h04;
im[1503]= 8'hCE;
im[1504]= 8'h93;
im[1505]= 8'h05;
im[1506]= 8'h04;
im[1507]= 8'hCD;
im[1508]= 8'h13;
im[1509]= 8'h06;
im[1510]= 8'h04;
im[1511]= 8'hCC;
im[1512]= 8'h03;
im[1513]= 8'h25;
im[1514]= 8'h04;
im[1515]= 8'hCE;
im[1516]= 8'h83;
im[1517]= 8'h25;
im[1518]= 8'h44;
im[1519]= 8'hCE;
im[1520]= 8'h03;
im[1521]= 8'h26;
im[1522]= 8'h84;
im[1523]= 8'hCE;
im[1524]= 8'h83;
im[1525]= 8'h26;
im[1526]= 8'hC4;
im[1527]= 8'hCE;
im[1528]= 8'h23;
im[1529]= 8'h2E;
im[1530]= 8'hD4;
im[1531]= 8'hF6;
im[1532]= 8'h23;
im[1533]= 8'h2C;
im[1534]= 8'hC4;
im[1535]= 8'hF6;
im[1536]= 8'h23;
im[1537]= 8'h2A;
im[1538]= 8'hB4;
im[1539]= 8'hF6;
im[1540]= 8'h23;
im[1541]= 8'h28;
im[1542]= 8'hA4;
im[1543]= 8'hF6;
im[1544]= 8'h03;
im[1545]= 8'h25;
im[1546]= 8'h04;
im[1547]= 8'hF7;
im[1548]= 8'h83;
im[1549]= 8'h25;
im[1550]= 8'h44;
im[1551]= 8'hF7;
im[1552]= 8'h03;
im[1553]= 8'h26;
im[1554]= 8'h84;
im[1555]= 8'hF7;
im[1556]= 8'h83;
im[1557]= 8'h26;
im[1558]= 8'hC4;
im[1559]= 8'hF7;
im[1560]= 8'h23;
im[1561]= 8'h2E;
im[1562]= 8'hD4;
im[1563]= 8'hC8;
im[1564]= 8'h23;
im[1565]= 8'h2C;
im[1566]= 8'hC4;
im[1567]= 8'hC8;
im[1568]= 8'h23;
im[1569]= 8'h2A;
im[1570]= 8'hB4;
im[1571]= 8'hC8;
im[1572]= 8'h23;
im[1573]= 8'h28;
im[1574]= 8'hA4;
im[1575]= 8'hC8;
im[1576]= 8'h23;
im[1577]= 8'h26;
im[1578]= 8'hD4;
im[1579]= 8'hCA;
im[1580]= 8'h23;
im[1581]= 8'h24;
im[1582]= 8'hC4;
im[1583]= 8'hCA;
im[1584]= 8'h23;
im[1585]= 8'h22;
im[1586]= 8'hB4;
im[1587]= 8'hCA;
im[1588]= 8'h23;
im[1589]= 8'h20;
im[1590]= 8'hA4;
im[1591]= 8'hCA;
im[1592]= 8'h13;
im[1593]= 8'h05;
im[1594]= 8'h04;
im[1595]= 8'hCB;
im[1596]= 8'h93;
im[1597]= 8'h05;
im[1598]= 8'h04;
im[1599]= 8'hCA;
im[1600]= 8'h13;
im[1601]= 8'h06;
im[1602]= 8'h04;
im[1603]= 8'hC9;
im[1604]= 8'h03;
im[1605]= 8'h25;
im[1606]= 8'h04;
im[1607]= 8'hCB;
im[1608]= 8'h23;
im[1609]= 8'h26;
im[1610]= 8'hA4;
im[1611]= 8'h84;
im[1612]= 8'h03;
im[1613]= 8'h25;
im[1614]= 8'h44;
im[1615]= 8'hCB;
im[1616]= 8'h23;
im[1617]= 8'h24;
im[1618]= 8'hA4;
im[1619]= 8'h84;
im[1620]= 8'h03;
im[1621]= 8'h25;
im[1622]= 8'h84;
im[1623]= 8'hCB;
im[1624]= 8'h23;
im[1625]= 8'h22;
im[1626]= 8'hA4;
im[1627]= 8'h84;
im[1628]= 8'h03;
im[1629]= 8'h25;
im[1630]= 8'hC4;
im[1631]= 8'hCB;
im[1632]= 8'h23;
im[1633]= 8'h20;
im[1634]= 8'hA4;
im[1635]= 8'h84;
im[1636]= 8'h03;
im[1637]= 8'h25;
im[1638]= 8'h04;
im[1639]= 8'hF8;
im[1640]= 8'h23;
im[1641]= 8'h2E;
im[1642]= 8'hA4;
im[1643]= 8'h82;
im[1644]= 8'h83;
im[1645]= 8'h25;
im[1646]= 8'h44;
im[1647]= 8'hF8;
im[1648]= 8'h23;
im[1649]= 8'h2C;
im[1650]= 8'hB4;
im[1651]= 8'h82;
im[1652]= 8'h03;
im[1653]= 8'h26;
im[1654]= 8'h84;
im[1655]= 8'hF8;
im[1656]= 8'h23;
im[1657]= 8'h2A;
im[1658]= 8'hC4;
im[1659]= 8'h82;
im[1660]= 8'h83;
im[1661]= 8'h26;
im[1662]= 8'hC4;
im[1663]= 8'hF8;
im[1664]= 8'h23;
im[1665]= 8'h28;
im[1666]= 8'hD4;
im[1667]= 8'h82;
im[1668]= 8'h23;
im[1669]= 8'h26;
im[1670]= 8'hD4;
im[1671]= 8'hC6;
im[1672]= 8'h23;
im[1673]= 8'h24;
im[1674]= 8'hC4;
im[1675]= 8'hC6;
im[1676]= 8'h23;
im[1677]= 8'h22;
im[1678]= 8'hB4;
im[1679]= 8'hC6;
im[1680]= 8'h23;
im[1681]= 8'h20;
im[1682]= 8'hA4;
im[1683]= 8'hC6;
im[1684]= 8'h23;
im[1685]= 8'h2E;
im[1686]= 8'hD4;
im[1687]= 8'hC6;
im[1688]= 8'h23;
im[1689]= 8'h2C;
im[1690]= 8'hC4;
im[1691]= 8'hC6;
im[1692]= 8'h23;
im[1693]= 8'h2A;
im[1694]= 8'hB4;
im[1695]= 8'hC6;
im[1696]= 8'h23;
im[1697]= 8'h28;
im[1698]= 8'hA4;
im[1699]= 8'hC6;
im[1700]= 8'h13;
im[1701]= 8'h05;
im[1702]= 8'h04;
im[1703]= 8'hC8;
im[1704]= 8'h93;
im[1705]= 8'h05;
im[1706]= 8'h04;
im[1707]= 8'hC7;
im[1708]= 8'h13;
im[1709]= 8'h06;
im[1710]= 8'h04;
im[1711]= 8'hC6;
im[1712]= 8'h83;
im[1713]= 8'h28;
im[1714]= 8'h04;
im[1715]= 8'h83;
im[1716]= 8'h03;
im[1717]= 8'h28;
im[1718]= 8'h44;
im[1719]= 8'h83;
im[1720]= 8'h83;
im[1721]= 8'h27;
im[1722]= 8'h84;
im[1723]= 8'h83;
im[1724]= 8'h03;
im[1725]= 8'h27;
im[1726]= 8'hC4;
im[1727]= 8'h83;
im[1728]= 8'h03;
im[1729]= 8'h25;
im[1730]= 8'h04;
im[1731]= 8'hC8;
im[1732]= 8'h83;
im[1733]= 8'h25;
im[1734]= 8'h44;
im[1735]= 8'hC8;
im[1736]= 8'h03;
im[1737]= 8'h26;
im[1738]= 8'h84;
im[1739]= 8'hC8;
im[1740]= 8'h83;
im[1741]= 8'h26;
im[1742]= 8'hC4;
im[1743]= 8'hC8;
im[1744]= 8'h23;
im[1745]= 8'h2E;
im[1746]= 8'h14;
im[1747]= 8'hC3;
im[1748]= 8'h23;
im[1749]= 8'h2C;
im[1750]= 8'h04;
im[1751]= 8'hC3;
im[1752]= 8'h23;
im[1753]= 8'h2A;
im[1754]= 8'hF4;
im[1755]= 8'hC2;
im[1756]= 8'h23;
im[1757]= 8'h28;
im[1758]= 8'hE4;
im[1759]= 8'hC2;
im[1760]= 8'h23;
im[1761]= 8'h26;
im[1762]= 8'hD4;
im[1763]= 8'hC4;
im[1764]= 8'h23;
im[1765]= 8'h24;
im[1766]= 8'hC4;
im[1767]= 8'hC4;
im[1768]= 8'h23;
im[1769]= 8'h22;
im[1770]= 8'hB4;
im[1771]= 8'hC4;
im[1772]= 8'h23;
im[1773]= 8'h20;
im[1774]= 8'hA4;
im[1775]= 8'hC4;
im[1776]= 8'h13;
im[1777]= 8'h05;
im[1778]= 8'h04;
im[1779]= 8'hC5;
im[1780]= 8'h93;
im[1781]= 8'h05;
im[1782]= 8'h04;
im[1783]= 8'hC4;
im[1784]= 8'h13;
im[1785]= 8'h06;
im[1786]= 8'h04;
im[1787]= 8'hC3;
im[1788]= 8'h83;
im[1789]= 8'h28;
im[1790]= 8'h04;
im[1791]= 8'h84;
im[1792]= 8'h03;
im[1793]= 8'h28;
im[1794]= 8'h44;
im[1795]= 8'h84;
im[1796]= 8'h83;
im[1797]= 8'h27;
im[1798]= 8'h84;
im[1799]= 8'h84;
im[1800]= 8'h03;
im[1801]= 8'h27;
im[1802]= 8'hC4;
im[1803]= 8'h84;
im[1804]= 8'h03;
im[1805]= 8'h25;
im[1806]= 8'h04;
im[1807]= 8'hC5;
im[1808]= 8'h83;
im[1809]= 8'h25;
im[1810]= 8'h44;
im[1811]= 8'hC5;
im[1812]= 8'h03;
im[1813]= 8'h26;
im[1814]= 8'h84;
im[1815]= 8'hC5;
im[1816]= 8'h83;
im[1817]= 8'h26;
im[1818]= 8'hC4;
im[1819]= 8'hC5;
im[1820]= 8'h23;
im[1821]= 8'h2E;
im[1822]= 8'h14;
im[1823]= 8'hC1;
im[1824]= 8'h23;
im[1825]= 8'h2C;
im[1826]= 8'h04;
im[1827]= 8'hC1;
im[1828]= 8'h23;
im[1829]= 8'h2A;
im[1830]= 8'hF4;
im[1831]= 8'hC0;
im[1832]= 8'h23;
im[1833]= 8'h28;
im[1834]= 8'hE4;
im[1835]= 8'hC0;
im[1836]= 8'h23;
im[1837]= 8'h26;
im[1838]= 8'hD4;
im[1839]= 8'hC0;
im[1840]= 8'h23;
im[1841]= 8'h24;
im[1842]= 8'hC4;
im[1843]= 8'hC0;
im[1844]= 8'h23;
im[1845]= 8'h22;
im[1846]= 8'hB4;
im[1847]= 8'hC0;
im[1848]= 8'h23;
im[1849]= 8'h20;
im[1850]= 8'hA4;
im[1851]= 8'hC0;
im[1852]= 8'h13;
im[1853]= 8'h05;
im[1854]= 8'h04;
im[1855]= 8'hC2;
im[1856]= 8'h93;
im[1857]= 8'h05;
im[1858]= 8'h04;
im[1859]= 8'hC1;
im[1860]= 8'h13;
im[1861]= 8'h06;
im[1862]= 8'h04;
im[1863]= 8'hC0;
im[1864]= 8'h03;
im[1865]= 8'h25;
im[1866]= 8'h04;
im[1867]= 8'hC2;
im[1868]= 8'h83;
im[1869]= 8'h25;
im[1870]= 8'h44;
im[1871]= 8'hC2;
im[1872]= 8'h03;
im[1873]= 8'h26;
im[1874]= 8'h84;
im[1875]= 8'hC2;
im[1876]= 8'h83;
im[1877]= 8'h26;
im[1878]= 8'hC4;
im[1879]= 8'hC2;
im[1880]= 8'h23;
im[1881]= 8'h2E;
im[1882]= 8'hD4;
im[1883]= 8'hBE;
im[1884]= 8'h23;
im[1885]= 8'h2C;
im[1886]= 8'hC4;
im[1887]= 8'hBE;
im[1888]= 8'h23;
im[1889]= 8'h2A;
im[1890]= 8'hB4;
im[1891]= 8'hBE;
im[1892]= 8'h23;
im[1893]= 8'h28;
im[1894]= 8'hA4;
im[1895]= 8'hBE;
im[1896]= 8'h13;
im[1897]= 8'h05;
im[1898]= 8'h04;
im[1899]= 8'hBF;
im[1900]= 8'h6F;
im[1901]= 8'h00;
im[1902]= 8'h40;
im[1903]= 8'h00;
im[1904]= 8'h83;
im[1905]= 8'h25;
im[1906]= 8'hC4;
im[1907]= 8'hFC;
im[1908]= 8'h13;
im[1909]= 8'h05;
im[1910]= 8'h30;
im[1911]= 8'h00;
im[1912]= 8'h23;
im[1913]= 8'hA0;
im[1914]= 8'hA5;
im[1915]= 8'h00;
im[1916]= 8'h03;
im[1917]= 8'h25;
im[1918]= 8'h04;
im[1919]= 8'hF7;
im[1920]= 8'h93;
im[1921]= 8'h85;
im[1922]= 8'h45;
im[1923]= 8'h76;
im[1924]= 8'hB3;
im[1925]= 8'h85;
im[1926]= 8'h85;
im[1927]= 8'h00;
im[1928]= 8'h23;
im[1929]= 8'hA0;
im[1930]= 8'hA5;
im[1931]= 8'h00;
im[1932]= 8'h03;
im[1933]= 8'h25;
im[1934]= 8'h44;
im[1935]= 8'hF7;
im[1936]= 8'h93;
im[1937]= 8'h85;
im[1938]= 8'h05;
im[1939]= 8'h76;
im[1940]= 8'hB3;
im[1941]= 8'h85;
im[1942]= 8'h85;
im[1943]= 8'h00;
im[1944]= 8'h23;
im[1945]= 8'hA0;
im[1946]= 8'hA5;
im[1947]= 8'h00;
im[1948]= 8'h03;
im[1949]= 8'h25;
im[1950]= 8'h84;
im[1951]= 8'hF7;
im[1952]= 8'h93;
im[1953]= 8'h85;
im[1954]= 8'hC5;
im[1955]= 8'h75;
im[1956]= 8'hB3;
im[1957]= 8'h85;
im[1958]= 8'h85;
im[1959]= 8'h00;
im[1960]= 8'h23;
im[1961]= 8'hA0;
im[1962]= 8'hA5;
im[1963]= 8'h00;
im[1964]= 8'h03;
im[1965]= 8'h25;
im[1966]= 8'hC4;
im[1967]= 8'hF7;
im[1968]= 8'h93;
im[1969]= 8'h85;
im[1970]= 8'h85;
im[1971]= 8'h75;
im[1972]= 8'hB3;
im[1973]= 8'h85;
im[1974]= 8'h85;
im[1975]= 8'h00;
im[1976]= 8'h23;
im[1977]= 8'hA0;
im[1978]= 8'hA5;
im[1979]= 8'h00;
im[1980]= 8'h03;
im[1981]= 8'h25;
im[1982]= 8'h04;
im[1983]= 8'hF8;
im[1984]= 8'h93;
im[1985]= 8'h85;
im[1986]= 8'h45;
im[1987]= 8'h75;
im[1988]= 8'hB3;
im[1989]= 8'h85;
im[1990]= 8'h85;
im[1991]= 8'h00;
im[1992]= 8'h23;
im[1993]= 8'hA0;
im[1994]= 8'hA5;
im[1995]= 8'h00;
im[1996]= 8'h83;
im[1997]= 8'h25;
im[1998]= 8'h44;
im[1999]= 8'hF8;
im[2000]= 8'h13;
im[2001]= 8'h06;
im[2002]= 8'h06;
im[2003]= 8'h75;
im[2004]= 8'h33;
im[2005]= 8'h06;
im[2006]= 8'h86;
im[2007]= 8'h00;
im[2008]= 8'h23;
im[2009]= 8'h20;
im[2010]= 8'hB6;
im[2011]= 8'h00;
im[2012]= 8'h03;
im[2013]= 8'h26;
im[2014]= 8'h84;
im[2015]= 8'hF8;
im[2016]= 8'h93;
im[2017]= 8'h86;
im[2018]= 8'hC6;
im[2019]= 8'h74;
im[2020]= 8'hB3;
im[2021]= 8'h86;
im[2022]= 8'h86;
im[2023]= 8'h00;
im[2024]= 8'h23;
im[2025]= 8'hA0;
im[2026]= 8'hC6;
im[2027]= 8'h00;
im[2028]= 8'h83;
im[2029]= 8'h26;
im[2030]= 8'hC4;
im[2031]= 8'hF8;
im[2032]= 8'h13;
im[2033]= 8'h07;
im[2034]= 8'h87;
im[2035]= 8'h74;
im[2036]= 8'h33;
im[2037]= 8'h07;
im[2038]= 8'h87;
im[2039]= 8'h00;
im[2040]= 8'h23;
im[2041]= 8'h20;
im[2042]= 8'hD7;
im[2043]= 8'h00;
im[2044]= 8'h23;
im[2045]= 8'h2E;
im[2046]= 8'hD4;
im[2047]= 8'hA6;
im[2048]= 8'h23;
im[2049]= 8'h2C;
im[2050]= 8'hC4;
im[2051]= 8'hA6;
im[2052]= 8'h23;
im[2053]= 8'h2A;
im[2054]= 8'hB4;
im[2055]= 8'hA6;
im[2056]= 8'h23;
im[2057]= 8'h28;
im[2058]= 8'hA4;
im[2059]= 8'hA6;
im[2060]= 8'h23;
im[2061]= 8'h26;
im[2062]= 8'hD4;
im[2063]= 8'hA8;
im[2064]= 8'h23;
im[2065]= 8'h24;
im[2066]= 8'hC4;
im[2067]= 8'hA8;
im[2068]= 8'h23;
im[2069]= 8'h22;
im[2070]= 8'hB4;
im[2071]= 8'hA8;
im[2072]= 8'h23;
im[2073]= 8'h20;
im[2074]= 8'hA4;
im[2075]= 8'hA8;
im[2076]= 8'h13;
im[2077]= 8'h05;
im[2078]= 8'h04;
im[2079]= 8'hA9;
im[2080]= 8'h93;
im[2081]= 8'h05;
im[2082]= 8'h04;
im[2083]= 8'hA8;
im[2084]= 8'h13;
im[2085]= 8'h06;
im[2086]= 8'h04;
im[2087]= 8'hA7;
im[2088]= 8'h13;
im[2089]= 8'h05;
im[2090]= 8'h85;
im[2091]= 8'h74;
im[2092]= 8'h33;
im[2093]= 8'h05;
im[2094]= 8'h85;
im[2095]= 8'h00;
im[2096]= 8'h83;
im[2097]= 8'h28;
im[2098]= 8'h05;
im[2099]= 8'h00;
im[2100]= 8'h13;
im[2101]= 8'h05;
im[2102]= 8'hC5;
im[2103]= 8'h74;
im[2104]= 8'h33;
im[2105]= 8'h05;
im[2106]= 8'h85;
im[2107]= 8'h00;
im[2108]= 8'h03;
im[2109]= 8'h28;
im[2110]= 8'h05;
im[2111]= 8'h00;
im[2112]= 8'h13;
im[2113]= 8'h05;
im[2114]= 8'h05;
im[2115]= 8'h75;
im[2116]= 8'h33;
im[2117]= 8'h05;
im[2118]= 8'h85;
im[2119]= 8'h00;
im[2120]= 8'h83;
im[2121]= 8'h27;
im[2122]= 8'h05;
im[2123]= 8'h00;
im[2124]= 8'h13;
im[2125]= 8'h05;
im[2126]= 8'h45;
im[2127]= 8'h75;
im[2128]= 8'h33;
im[2129]= 8'h05;
im[2130]= 8'h85;
im[2131]= 8'h00;
im[2132]= 8'h03;
im[2133]= 8'h27;
im[2134]= 8'h05;
im[2135]= 8'h00;
im[2136]= 8'h03;
im[2137]= 8'h25;
im[2138]= 8'h04;
im[2139]= 8'hA9;
im[2140]= 8'h83;
im[2141]= 8'h25;
im[2142]= 8'h44;
im[2143]= 8'hA9;
im[2144]= 8'h03;
im[2145]= 8'h26;
im[2146]= 8'h84;
im[2147]= 8'hA9;
im[2148]= 8'h83;
im[2149]= 8'h26;
im[2150]= 8'hC4;
im[2151]= 8'hA9;
im[2152]= 8'h23;
im[2153]= 8'h26;
im[2154]= 8'h14;
im[2155]= 8'hA5;
im[2156]= 8'h23;
im[2157]= 8'h24;
im[2158]= 8'h04;
im[2159]= 8'hA5;
im[2160]= 8'h23;
im[2161]= 8'h22;
im[2162]= 8'hF4;
im[2163]= 8'hA4;
im[2164]= 8'h23;
im[2165]= 8'h20;
im[2166]= 8'hE4;
im[2167]= 8'hA4;
im[2168]= 8'h23;
im[2169]= 8'h2E;
im[2170]= 8'hD4;
im[2171]= 8'hA4;
im[2172]= 8'h23;
im[2173]= 8'h2C;
im[2174]= 8'hC4;
im[2175]= 8'hA4;
im[2176]= 8'h23;
im[2177]= 8'h2A;
im[2178]= 8'hB4;
im[2179]= 8'hA4;
im[2180]= 8'h23;
im[2181]= 8'h28;
im[2182]= 8'hA4;
im[2183]= 8'hA4;
im[2184]= 8'h13;
im[2185]= 8'h05;
im[2186]= 8'h04;
im[2187]= 8'hA6;
im[2188]= 8'h93;
im[2189]= 8'h05;
im[2190]= 8'h04;
im[2191]= 8'hA5;
im[2192]= 8'h13;
im[2193]= 8'h06;
im[2194]= 8'h04;
im[2195]= 8'hA4;
im[2196]= 8'h03;
im[2197]= 8'h25;
im[2198]= 8'h04;
im[2199]= 8'hA6;
im[2200]= 8'h83;
im[2201]= 8'h25;
im[2202]= 8'h44;
im[2203]= 8'hA6;
im[2204]= 8'h03;
im[2205]= 8'h26;
im[2206]= 8'h84;
im[2207]= 8'hA6;
im[2208]= 8'h83;
im[2209]= 8'h26;
im[2210]= 8'hC4;
im[2211]= 8'hA6;
im[2212]= 8'h23;
im[2213]= 8'h26;
im[2214]= 8'hD4;
im[2215]= 8'hAA;
im[2216]= 8'h23;
im[2217]= 8'h24;
im[2218]= 8'hC4;
im[2219]= 8'hAA;
im[2220]= 8'h23;
im[2221]= 8'h22;
im[2222]= 8'hB4;
im[2223]= 8'hAA;
im[2224]= 8'h23;
im[2225]= 8'h20;
im[2226]= 8'hA4;
im[2227]= 8'hAA;
im[2228]= 8'h13;
im[2229]= 8'h05;
im[2230]= 8'h04;
im[2231]= 8'hAB;
im[2232]= 8'h93;
im[2233]= 8'h05;
im[2234]= 8'h04;
im[2235]= 8'hAA;
im[2236]= 8'h13;
im[2237]= 8'h05;
im[2238]= 8'h85;
im[2239]= 8'h75;
im[2240]= 8'h33;
im[2241]= 8'h05;
im[2242]= 8'h85;
im[2243]= 8'h00;
im[2244]= 8'h83;
im[2245]= 8'h28;
im[2246]= 8'h05;
im[2247]= 8'h00;
im[2248]= 8'h13;
im[2249]= 8'h05;
im[2250]= 8'hC5;
im[2251]= 8'h75;
im[2252]= 8'h33;
im[2253]= 8'h05;
im[2254]= 8'h85;
im[2255]= 8'h00;
im[2256]= 8'h03;
im[2257]= 8'h28;
im[2258]= 8'h05;
im[2259]= 8'h00;
im[2260]= 8'h13;
im[2261]= 8'h05;
im[2262]= 8'h05;
im[2263]= 8'h76;
im[2264]= 8'h33;
im[2265]= 8'h05;
im[2266]= 8'h85;
im[2267]= 8'h00;
im[2268]= 8'h83;
im[2269]= 8'h27;
im[2270]= 8'h05;
im[2271]= 8'h00;
im[2272]= 8'h13;
im[2273]= 8'h05;
im[2274]= 8'h45;
im[2275]= 8'h76;
im[2276]= 8'h33;
im[2277]= 8'h05;
im[2278]= 8'h85;
im[2279]= 8'h00;
im[2280]= 8'h03;
im[2281]= 8'h27;
im[2282]= 8'h05;
im[2283]= 8'h00;
im[2284]= 8'h03;
im[2285]= 8'h25;
im[2286]= 8'h04;
im[2287]= 8'hAB;
im[2288]= 8'h83;
im[2289]= 8'h25;
im[2290]= 8'h44;
im[2291]= 8'hAB;
im[2292]= 8'h03;
im[2293]= 8'h26;
im[2294]= 8'h84;
im[2295]= 8'hAB;
im[2296]= 8'h83;
im[2297]= 8'h26;
im[2298]= 8'hC4;
im[2299]= 8'hAB;
im[2300]= 8'h23;
im[2301]= 8'h26;
im[2302]= 8'h14;
im[2303]= 8'hA3;
im[2304]= 8'h23;
im[2305]= 8'h24;
im[2306]= 8'h04;
im[2307]= 8'hA3;
im[2308]= 8'h23;
im[2309]= 8'h22;
im[2310]= 8'hF4;
im[2311]= 8'hA2;
im[2312]= 8'h23;
im[2313]= 8'h20;
im[2314]= 8'hE4;
im[2315]= 8'hA2;
im[2316]= 8'h23;
im[2317]= 8'h2E;
im[2318]= 8'hD4;
im[2319]= 8'hA0;
im[2320]= 8'h23;
im[2321]= 8'h2C;
im[2322]= 8'hC4;
im[2323]= 8'hA0;
im[2324]= 8'h23;
im[2325]= 8'h2A;
im[2326]= 8'hB4;
im[2327]= 8'hA0;
im[2328]= 8'h23;
im[2329]= 8'h28;
im[2330]= 8'hA4;
im[2331]= 8'hA0;
im[2332]= 8'h13;
im[2333]= 8'h05;
im[2334]= 8'h04;
im[2335]= 8'hA3;
im[2336]= 8'h93;
im[2337]= 8'h05;
im[2338]= 8'h04;
im[2339]= 8'hA2;
im[2340]= 8'h13;
im[2341]= 8'h06;
im[2342]= 8'h04;
im[2343]= 8'hA1;
im[2344]= 8'h03;
im[2345]= 8'h25;
im[2346]= 8'h04;
im[2347]= 8'hA3;
im[2348]= 8'h83;
im[2349]= 8'h25;
im[2350]= 8'h44;
im[2351]= 8'hA3;
im[2352]= 8'h03;
im[2353]= 8'h26;
im[2354]= 8'h84;
im[2355]= 8'hA3;
im[2356]= 8'h83;
im[2357]= 8'h26;
im[2358]= 8'hC4;
im[2359]= 8'hA3;
im[2360]= 8'h23;
im[2361]= 8'h26;
im[2362]= 8'hD4;
im[2363]= 8'hA0;
im[2364]= 8'h23;
im[2365]= 8'h24;
im[2366]= 8'hC4;
im[2367]= 8'hA0;
im[2368]= 8'h23;
im[2369]= 8'h22;
im[2370]= 8'hB4;
im[2371]= 8'hA0;
im[2372]= 8'h23;
im[2373]= 8'h20;
im[2374]= 8'hA4;
im[2375]= 8'hA0;
im[2376]= 8'h13;
im[2377]= 8'h05;
im[2378]= 8'h04;
im[2379]= 8'hA0;
im[2380]= 8'h03;
im[2381]= 8'h25;
im[2382]= 8'h04;
im[2383]= 8'hF8;
im[2384]= 8'h83;
im[2385]= 8'h25;
im[2386]= 8'h44;
im[2387]= 8'hF8;
im[2388]= 8'h03;
im[2389]= 8'h26;
im[2390]= 8'h84;
im[2391]= 8'hF8;
im[2392]= 8'h83;
im[2393]= 8'h26;
im[2394]= 8'hC4;
im[2395]= 8'hF8;
im[2396]= 8'h23;
im[2397]= 8'h2E;
im[2398]= 8'hD4;
im[2399]= 8'h9E;
im[2400]= 8'h23;
im[2401]= 8'h2C;
im[2402]= 8'hC4;
im[2403]= 8'h9E;
im[2404]= 8'h23;
im[2405]= 8'h2A;
im[2406]= 8'hB4;
im[2407]= 8'h9E;
im[2408]= 8'h23;
im[2409]= 8'h28;
im[2410]= 8'hA4;
im[2411]= 8'h9E;
im[2412]= 8'h13;
im[2413]= 8'h05;
im[2414]= 8'h04;
im[2415]= 8'h9F;
im[2416]= 8'h13;
im[2417]= 8'h05;
im[2418]= 8'h05;
im[2419]= 8'h7A;
im[2420]= 8'h33;
im[2421]= 8'h05;
im[2422]= 8'h85;
im[2423]= 8'h00;
im[2424]= 8'h13;
im[2425]= 8'h05;
im[2426]= 8'h85;
im[2427]= 8'h76;
im[2428]= 8'h33;
im[2429]= 8'h05;
im[2430]= 8'h85;
im[2431]= 8'h00;
im[2432]= 8'h13;
im[2433]= 8'h05;
im[2434]= 8'h05;
im[2435]= 8'h7C;
im[2436]= 8'h33;
im[2437]= 8'h05;
im[2438]= 8'h85;
im[2439]= 8'h00;
im[2440]= 8'h13;
im[2441]= 8'h05;
im[2442]= 8'h85;
im[2443]= 8'h76;
im[2444]= 8'h33;
im[2445]= 8'h05;
im[2446]= 8'h85;
im[2447]= 8'h00;
im[2448]= 8'h13;
im[2449]= 8'h05;
im[2450]= 8'h04;
im[2451]= 8'h9E;
im[2452]= 8'h03;
im[2453]= 8'h25;
im[2454]= 8'h04;
im[2455]= 8'h9E;
im[2456]= 8'h93;
im[2457]= 8'h85;
im[2458]= 8'hC5;
im[2459]= 8'h77;
im[2460]= 8'hB3;
im[2461]= 8'h85;
im[2462]= 8'h85;
im[2463]= 8'h00;
im[2464]= 8'h23;
im[2465]= 8'hA0;
im[2466]= 8'hA5;
im[2467]= 8'h00;
im[2468]= 8'h03;
im[2469]= 8'h25;
im[2470]= 8'h44;
im[2471]= 8'h9E;
im[2472]= 8'h93;
im[2473]= 8'h85;
im[2474]= 8'h85;
im[2475]= 8'h77;
im[2476]= 8'hB3;
im[2477]= 8'h85;
im[2478]= 8'h85;
im[2479]= 8'h00;
im[2480]= 8'h23;
im[2481]= 8'hA0;
im[2482]= 8'hA5;
im[2483]= 8'h00;
im[2484]= 8'h03;
im[2485]= 8'h25;
im[2486]= 8'h84;
im[2487]= 8'h9E;
im[2488]= 8'h93;
im[2489]= 8'h85;
im[2490]= 8'h45;
im[2491]= 8'h77;
im[2492]= 8'hB3;
im[2493]= 8'h85;
im[2494]= 8'h85;
im[2495]= 8'h00;
im[2496]= 8'h23;
im[2497]= 8'hA0;
im[2498]= 8'hA5;
im[2499]= 8'h00;
im[2500]= 8'h03;
im[2501]= 8'h25;
im[2502]= 8'hC4;
im[2503]= 8'h9E;
im[2504]= 8'h93;
im[2505]= 8'h85;
im[2506]= 8'h05;
im[2507]= 8'h77;
im[2508]= 8'hB3;
im[2509]= 8'h85;
im[2510]= 8'h85;
im[2511]= 8'h00;
im[2512]= 8'h23;
im[2513]= 8'hA0;
im[2514]= 8'hA5;
im[2515]= 8'h00;
im[2516]= 8'h03;
im[2517]= 8'h25;
im[2518]= 8'h04;
im[2519]= 8'hFB;
im[2520]= 8'h83;
im[2521]= 8'h25;
im[2522]= 8'h44;
im[2523]= 8'hFB;
im[2524]= 8'h03;
im[2525]= 8'h26;
im[2526]= 8'h84;
im[2527]= 8'hFB;
im[2528]= 8'h83;
im[2529]= 8'h26;
im[2530]= 8'hC4;
im[2531]= 8'hFB;
im[2532]= 8'h93;
im[2533]= 8'h87;
im[2534]= 8'h07;
im[2535]= 8'h7D;
im[2536]= 8'hB3;
im[2537]= 8'h87;
im[2538]= 8'h87;
im[2539]= 8'h00;
im[2540]= 8'h23;
im[2541]= 8'hA0;
im[2542]= 8'hE7;
im[2543]= 8'h00;
im[2544]= 8'h23;
im[2545]= 8'h2E;
im[2546]= 8'hE4;
im[2547]= 8'h9A;
im[2548]= 8'h93;
im[2549]= 8'h87;
im[2550]= 8'h47;
im[2551]= 8'h7D;
im[2552]= 8'hB3;
im[2553]= 8'h87;
im[2554]= 8'h87;
im[2555]= 8'h00;
im[2556]= 8'h23;
im[2557]= 8'hA0;
im[2558]= 8'hE7;
im[2559]= 8'h00;
im[2560]= 8'h23;
im[2561]= 8'h2C;
im[2562]= 8'hE4;
im[2563]= 8'h9A;
im[2564]= 8'h23;
im[2565]= 8'h2A;
im[2566]= 8'hE4;
im[2567]= 8'h9A;
im[2568]= 8'h23;
im[2569]= 8'h28;
im[2570]= 8'hE4;
im[2571]= 8'h9A;
im[2572]= 8'h23;
im[2573]= 8'h26;
im[2574]= 8'hD4;
im[2575]= 8'h9C;
im[2576]= 8'h23;
im[2577]= 8'h24;
im[2578]= 8'hC4;
im[2579]= 8'h9C;
im[2580]= 8'h23;
im[2581]= 8'h22;
im[2582]= 8'hB4;
im[2583]= 8'h9C;
im[2584]= 8'h23;
im[2585]= 8'h20;
im[2586]= 8'hA4;
im[2587]= 8'h9C;
im[2588]= 8'h13;
im[2589]= 8'h05;
im[2590]= 8'h04;
im[2591]= 8'h9D;
im[2592]= 8'h93;
im[2593]= 8'h05;
im[2594]= 8'h04;
im[2595]= 8'h9C;
im[2596]= 8'h13;
im[2597]= 8'h06;
im[2598]= 8'h04;
im[2599]= 8'h9B;
im[2600]= 8'h13;
im[2601]= 8'h05;
im[2602]= 8'h05;
im[2603]= 8'h77;
im[2604]= 8'h33;
im[2605]= 8'h05;
im[2606]= 8'h85;
im[2607]= 8'h00;
im[2608]= 8'h83;
im[2609]= 8'h28;
im[2610]= 8'h05;
im[2611]= 8'h00;
im[2612]= 8'h13;
im[2613]= 8'h05;
im[2614]= 8'h45;
im[2615]= 8'h77;
im[2616]= 8'h33;
im[2617]= 8'h05;
im[2618]= 8'h85;
im[2619]= 8'h00;
im[2620]= 8'h03;
im[2621]= 8'h28;
im[2622]= 8'h05;
im[2623]= 8'h00;
im[2624]= 8'h13;
im[2625]= 8'h05;
im[2626]= 8'h85;
im[2627]= 8'h77;
im[2628]= 8'h33;
im[2629]= 8'h05;
im[2630]= 8'h85;
im[2631]= 8'h00;
im[2632]= 8'h83;
im[2633]= 8'h27;
im[2634]= 8'h05;
im[2635]= 8'h00;
im[2636]= 8'h13;
im[2637]= 8'h05;
im[2638]= 8'hC5;
im[2639]= 8'h77;
im[2640]= 8'h33;
im[2641]= 8'h05;
im[2642]= 8'h85;
im[2643]= 8'h00;
im[2644]= 8'h03;
im[2645]= 8'h27;
im[2646]= 8'h05;
im[2647]= 8'h00;
im[2648]= 8'h03;
im[2649]= 8'h25;
im[2650]= 8'h04;
im[2651]= 8'h9D;
im[2652]= 8'h83;
im[2653]= 8'h25;
im[2654]= 8'h44;
im[2655]= 8'h9D;
im[2656]= 8'h03;
im[2657]= 8'h26;
im[2658]= 8'h84;
im[2659]= 8'h9D;
im[2660]= 8'h83;
im[2661]= 8'h26;
im[2662]= 8'hC4;
im[2663]= 8'h9D;
im[2664]= 8'h23;
im[2665]= 8'h2E;
im[2666]= 8'h14;
im[2667]= 8'h99;
im[2668]= 8'h23;
im[2669]= 8'h2C;
im[2670]= 8'h04;
im[2671]= 8'h99;
im[2672]= 8'h23;
im[2673]= 8'h2A;
im[2674]= 8'hF4;
im[2675]= 8'h98;
im[2676]= 8'h23;
im[2677]= 8'h28;
im[2678]= 8'hE4;
im[2679]= 8'h98;
im[2680]= 8'h23;
im[2681]= 8'h26;
im[2682]= 8'hD4;
im[2683]= 8'h98;
im[2684]= 8'h23;
im[2685]= 8'h24;
im[2686]= 8'hC4;
im[2687]= 8'h98;
im[2688]= 8'h23;
im[2689]= 8'h22;
im[2690]= 8'hB4;
im[2691]= 8'h98;
im[2692]= 8'h23;
im[2693]= 8'h20;
im[2694]= 8'hA4;
im[2695]= 8'h98;
im[2696]= 8'h13;
im[2697]= 8'h05;
im[2698]= 8'h04;
im[2699]= 8'h9A;
im[2700]= 8'h93;
im[2701]= 8'h05;
im[2702]= 8'h04;
im[2703]= 8'h99;
im[2704]= 8'h13;
im[2705]= 8'h06;
im[2706]= 8'h04;
im[2707]= 8'h98;
im[2708]= 8'h03;
im[2709]= 8'h25;
im[2710]= 8'h04;
im[2711]= 8'h9A;
im[2712]= 8'h83;
im[2713]= 8'h25;
im[2714]= 8'h44;
im[2715]= 8'h9A;
im[2716]= 8'h03;
im[2717]= 8'h26;
im[2718]= 8'h84;
im[2719]= 8'h9A;
im[2720]= 8'h83;
im[2721]= 8'h26;
im[2722]= 8'hC4;
im[2723]= 8'h9A;
im[2724]= 8'h23;
im[2725]= 8'h2E;
im[2726]= 8'hD4;
im[2727]= 8'h96;
im[2728]= 8'h23;
im[2729]= 8'h2C;
im[2730]= 8'hC4;
im[2731]= 8'h96;
im[2732]= 8'h23;
im[2733]= 8'h2A;
im[2734]= 8'hB4;
im[2735]= 8'h96;
im[2736]= 8'h23;
im[2737]= 8'h28;
im[2738]= 8'hA4;
im[2739]= 8'h96;
im[2740]= 8'h13;
im[2741]= 8'h05;
im[2742]= 8'h04;
im[2743]= 8'h97;
im[2744]= 8'h03;
im[2745]= 8'h25;
im[2746]= 8'h84;
im[2747]= 8'hFC;
im[2748]= 8'h03;
im[2749]= 8'h25;
im[2750]= 8'h04;
im[2751]= 8'hF8;
im[2752]= 8'h83;
im[2753]= 8'h25;
im[2754]= 8'h44;
im[2755]= 8'hF8;
im[2756]= 8'h03;
im[2757]= 8'h26;
im[2758]= 8'h84;
im[2759]= 8'hF8;
im[2760]= 8'h83;
im[2761]= 8'h26;
im[2762]= 8'hC4;
im[2763]= 8'hF8;
im[2764]= 8'h23;
im[2765]= 8'h26;
im[2766]= 8'hD4;
im[2767]= 8'h96;
im[2768]= 8'h23;
im[2769]= 8'h24;
im[2770]= 8'hC4;
im[2771]= 8'h96;
im[2772]= 8'h23;
im[2773]= 8'h22;
im[2774]= 8'hB4;
im[2775]= 8'h96;
im[2776]= 8'h23;
im[2777]= 8'h20;
im[2778]= 8'hA4;
im[2779]= 8'h96;
im[2780]= 8'h13;
im[2781]= 8'h05;
im[2782]= 8'h04;
im[2783]= 8'h96;
im[2784]= 8'h13;
im[2785]= 8'h05;
im[2786]= 8'h05;
im[2787]= 8'h7A;
im[2788]= 8'h33;
im[2789]= 8'h05;
im[2790]= 8'h85;
im[2791]= 8'h00;
im[2792]= 8'h13;
im[2793]= 8'h05;
im[2794]= 8'h85;
im[2795]= 8'h78;
im[2796]= 8'h33;
im[2797]= 8'h05;
im[2798]= 8'h85;
im[2799]= 8'h00;
im[2800]= 8'h13;
im[2801]= 8'h05;
im[2802]= 8'h05;
im[2803]= 8'h78;
im[2804]= 8'h33;
im[2805]= 8'h05;
im[2806]= 8'h85;
im[2807]= 8'h00;
im[2808]= 8'h13;
im[2809]= 8'h05;
im[2810]= 8'h85;
im[2811]= 8'h7A;
im[2812]= 8'h33;
im[2813]= 8'h05;
im[2814]= 8'h85;
im[2815]= 8'h00;
im[2816]= 8'h13;
im[2817]= 8'h05;
im[2818]= 8'h05;
im[2819]= 8'h78;
im[2820]= 8'h33;
im[2821]= 8'h05;
im[2822]= 8'h85;
im[2823]= 8'h00;
im[2824]= 8'h13;
im[2825]= 8'h05;
im[2826]= 8'h05;
im[2827]= 8'h7C;
im[2828]= 8'h33;
im[2829]= 8'h05;
im[2830]= 8'h85;
im[2831]= 8'h00;
im[2832]= 8'h13;
im[2833]= 8'h05;
im[2834]= 8'h05;
im[2835]= 8'h7B;
im[2836]= 8'h33;
im[2837]= 8'h05;
im[2838]= 8'h85;
im[2839]= 8'h00;
im[2840]= 8'h13;
im[2841]= 8'h05;
im[2842]= 8'h85;
im[2843]= 8'h78;
im[2844]= 8'h33;
im[2845]= 8'h05;
im[2846]= 8'h85;
im[2847]= 8'h00;
im[2848]= 8'h13;
im[2849]= 8'h05;
im[2850]= 8'h04;
im[2851]= 8'h95;
im[2852]= 8'h13;
im[2853]= 8'h05;
im[2854]= 8'h05;
im[2855]= 8'h7D;
im[2856]= 8'h33;
im[2857]= 8'h05;
im[2858]= 8'h85;
im[2859]= 8'h00;
im[2860]= 8'h83;
im[2861]= 8'h27;
im[2862]= 8'h05;
im[2863]= 8'h00;
im[2864]= 8'h13;
im[2865]= 8'h05;
im[2866]= 8'h45;
im[2867]= 8'h7D;
im[2868]= 8'h33;
im[2869]= 8'h05;
im[2870]= 8'h85;
im[2871]= 8'h00;
im[2872]= 8'h03;
im[2873]= 8'h27;
im[2874]= 8'h05;
im[2875]= 8'h00;
im[2876]= 8'h03;
im[2877]= 8'h25;
im[2878]= 8'h04;
im[2879]= 8'h95;
im[2880]= 8'h93;
im[2881]= 8'h85;
im[2882]= 8'hC5;
im[2883]= 8'h79;
im[2884]= 8'hB3;
im[2885]= 8'h85;
im[2886]= 8'h85;
im[2887]= 8'h00;
im[2888]= 8'h23;
im[2889]= 8'hA0;
im[2890]= 8'hA5;
im[2891]= 8'h00;
im[2892]= 8'h03;
im[2893]= 8'h25;
im[2894]= 8'h44;
im[2895]= 8'h95;
im[2896]= 8'h93;
im[2897]= 8'h85;
im[2898]= 8'h85;
im[2899]= 8'h79;
im[2900]= 8'hB3;
im[2901]= 8'h85;
im[2902]= 8'h85;
im[2903]= 8'h00;
im[2904]= 8'h23;
im[2905]= 8'hA0;
im[2906]= 8'hA5;
im[2907]= 8'h00;
im[2908]= 8'h03;
im[2909]= 8'h25;
im[2910]= 8'h84;
im[2911]= 8'h95;
im[2912]= 8'h93;
im[2913]= 8'h85;
im[2914]= 8'h45;
im[2915]= 8'h79;
im[2916]= 8'hB3;
im[2917]= 8'h85;
im[2918]= 8'h85;
im[2919]= 8'h00;
im[2920]= 8'h23;
im[2921]= 8'hA0;
im[2922]= 8'hA5;
im[2923]= 8'h00;
im[2924]= 8'h03;
im[2925]= 8'h25;
im[2926]= 8'hC4;
im[2927]= 8'h95;
im[2928]= 8'h93;
im[2929]= 8'h85;
im[2930]= 8'h05;
im[2931]= 8'h79;
im[2932]= 8'hB3;
im[2933]= 8'h85;
im[2934]= 8'h85;
im[2935]= 8'h00;
im[2936]= 8'h23;
im[2937]= 8'hA0;
im[2938]= 8'hA5;
im[2939]= 8'h00;
im[2940]= 8'h03;
im[2941]= 8'h25;
im[2942]= 8'h04;
im[2943]= 8'hFB;
im[2944]= 8'h83;
im[2945]= 8'h25;
im[2946]= 8'h44;
im[2947]= 8'hFB;
im[2948]= 8'h03;
im[2949]= 8'h26;
im[2950]= 8'h84;
im[2951]= 8'hFB;
im[2952]= 8'h83;
im[2953]= 8'h26;
im[2954]= 8'hC4;
im[2955]= 8'hFB;
im[2956]= 8'h23;
im[2957]= 8'h26;
im[2958]= 8'hF4;
im[2959]= 8'h92;
im[2960]= 8'h23;
im[2961]= 8'h24;
im[2962]= 8'hE4;
im[2963]= 8'h92;
im[2964]= 8'h23;
im[2965]= 8'h22;
im[2966]= 8'hE4;
im[2967]= 8'h92;
im[2968]= 8'h23;
im[2969]= 8'h20;
im[2970]= 8'hE4;
im[2971]= 8'h92;
im[2972]= 8'h23;
im[2973]= 8'h2E;
im[2974]= 8'hD4;
im[2975]= 8'h92;
im[2976]= 8'h23;
im[2977]= 8'h2C;
im[2978]= 8'hC4;
im[2979]= 8'h92;
im[2980]= 8'h23;
im[2981]= 8'h2A;
im[2982]= 8'hB4;
im[2983]= 8'h92;
im[2984]= 8'h23;
im[2985]= 8'h28;
im[2986]= 8'hA4;
im[2987]= 8'h92;
im[2988]= 8'h13;
im[2989]= 8'h05;
im[2990]= 8'h04;
im[2991]= 8'h94;
im[2992]= 8'h93;
im[2993]= 8'h05;
im[2994]= 8'h04;
im[2995]= 8'h93;
im[2996]= 8'h13;
im[2997]= 8'h06;
im[2998]= 8'h04;
im[2999]= 8'h92;
im[3000]= 8'h13;
im[3001]= 8'h05;
im[3002]= 8'h05;
im[3003]= 8'h79;
im[3004]= 8'h33;
im[3005]= 8'h05;
im[3006]= 8'h85;
im[3007]= 8'h00;
im[3008]= 8'h83;
im[3009]= 8'h28;
im[3010]= 8'h05;
im[3011]= 8'h00;
im[3012]= 8'h13;
im[3013]= 8'h05;
im[3014]= 8'h45;
im[3015]= 8'h79;
im[3016]= 8'h33;
im[3017]= 8'h05;
im[3018]= 8'h85;
im[3019]= 8'h00;
im[3020]= 8'h03;
im[3021]= 8'h28;
im[3022]= 8'h05;
im[3023]= 8'h00;
im[3024]= 8'h13;
im[3025]= 8'h05;
im[3026]= 8'h85;
im[3027]= 8'h79;
im[3028]= 8'h33;
im[3029]= 8'h05;
im[3030]= 8'h85;
im[3031]= 8'h00;
im[3032]= 8'h83;
im[3033]= 8'h27;
im[3034]= 8'h05;
im[3035]= 8'h00;
im[3036]= 8'h13;
im[3037]= 8'h05;
im[3038]= 8'hC5;
im[3039]= 8'h79;
im[3040]= 8'h33;
im[3041]= 8'h05;
im[3042]= 8'h85;
im[3043]= 8'h00;
im[3044]= 8'h03;
im[3045]= 8'h27;
im[3046]= 8'h05;
im[3047]= 8'h00;
im[3048]= 8'h03;
im[3049]= 8'h25;
im[3050]= 8'h04;
im[3051]= 8'h94;
im[3052]= 8'h83;
im[3053]= 8'h25;
im[3054]= 8'h44;
im[3055]= 8'h94;
im[3056]= 8'h03;
im[3057]= 8'h26;
im[3058]= 8'h84;
im[3059]= 8'h94;
im[3060]= 8'h83;
im[3061]= 8'h26;
im[3062]= 8'hC4;
im[3063]= 8'h94;
im[3064]= 8'h23;
im[3065]= 8'h26;
im[3066]= 8'h14;
im[3067]= 8'h91;
im[3068]= 8'h23;
im[3069]= 8'h24;
im[3070]= 8'h04;
im[3071]= 8'h91;
im[3072]= 8'h23;
im[3073]= 8'h22;
im[3074]= 8'hF4;
im[3075]= 8'h90;
im[3076]= 8'h23;
im[3077]= 8'h20;
im[3078]= 8'hE4;
im[3079]= 8'h90;
im[3080]= 8'h23;
im[3081]= 8'h2E;
im[3082]= 8'hD4;
im[3083]= 8'h8E;
im[3084]= 8'h23;
im[3085]= 8'h2C;
im[3086]= 8'hC4;
im[3087]= 8'h8E;
im[3088]= 8'h23;
im[3089]= 8'h2A;
im[3090]= 8'hB4;
im[3091]= 8'h8E;
im[3092]= 8'h23;
im[3093]= 8'h28;
im[3094]= 8'hA4;
im[3095]= 8'h8E;
im[3096]= 8'h13;
im[3097]= 8'h05;
im[3098]= 8'h04;
im[3099]= 8'h91;
im[3100]= 8'h93;
im[3101]= 8'h05;
im[3102]= 8'h04;
im[3103]= 8'h90;
im[3104]= 8'h13;
im[3105]= 8'h06;
im[3106]= 8'h04;
im[3107]= 8'h8F;
im[3108]= 8'h03;
im[3109]= 8'h25;
im[3110]= 8'h04;
im[3111]= 8'h91;
im[3112]= 8'h83;
im[3113]= 8'h25;
im[3114]= 8'h44;
im[3115]= 8'h91;
im[3116]= 8'h03;
im[3117]= 8'h26;
im[3118]= 8'h84;
im[3119]= 8'h91;
im[3120]= 8'h83;
im[3121]= 8'h26;
im[3122]= 8'hC4;
im[3123]= 8'h91;
im[3124]= 8'h23;
im[3125]= 8'h26;
im[3126]= 8'hD4;
im[3127]= 8'h8E;
im[3128]= 8'h23;
im[3129]= 8'h24;
im[3130]= 8'hC4;
im[3131]= 8'h8E;
im[3132]= 8'h23;
im[3133]= 8'h22;
im[3134]= 8'hB4;
im[3135]= 8'h8E;
im[3136]= 8'h23;
im[3137]= 8'h20;
im[3138]= 8'hA4;
im[3139]= 8'h8E;
im[3140]= 8'h13;
im[3141]= 8'h05;
im[3142]= 8'h04;
im[3143]= 8'h8E;
im[3144]= 8'h03;
im[3145]= 8'h25;
im[3146]= 8'h84;
im[3147]= 8'hFC;
im[3148]= 8'h03;
im[3149]= 8'h25;
im[3150]= 8'h04;
im[3151]= 8'hF8;
im[3152]= 8'h83;
im[3153]= 8'h25;
im[3154]= 8'h44;
im[3155]= 8'hF8;
im[3156]= 8'h03;
im[3157]= 8'h26;
im[3158]= 8'h84;
im[3159]= 8'hF8;
im[3160]= 8'h83;
im[3161]= 8'h26;
im[3162]= 8'hC4;
im[3163]= 8'hF8;
im[3164]= 8'h23;
im[3165]= 8'h2E;
im[3166]= 8'hD4;
im[3167]= 8'h8C;
im[3168]= 8'h23;
im[3169]= 8'h2C;
im[3170]= 8'hC4;
im[3171]= 8'h8C;
im[3172]= 8'h23;
im[3173]= 8'h2A;
im[3174]= 8'hB4;
im[3175]= 8'h8C;
im[3176]= 8'h23;
im[3177]= 8'h28;
im[3178]= 8'hA4;
im[3179]= 8'h8C;
im[3180]= 8'h13;
im[3181]= 8'h05;
im[3182]= 8'h04;
im[3183]= 8'h8D;
im[3184]= 8'h13;
im[3185]= 8'h05;
im[3186]= 8'h05;
im[3187]= 8'h7A;
im[3188]= 8'h33;
im[3189]= 8'h05;
im[3190]= 8'h85;
im[3191]= 8'h00;
im[3192]= 8'h13;
im[3193]= 8'h05;
im[3194]= 8'h85;
im[3195]= 8'h7A;
im[3196]= 8'h33;
im[3197]= 8'h05;
im[3198]= 8'h85;
im[3199]= 8'h00;
im[3200]= 8'h13;
im[3201]= 8'h05;
im[3202]= 8'h85;
im[3203]= 8'h7C;
im[3204]= 8'h33;
im[3205]= 8'h05;
im[3206]= 8'h85;
im[3207]= 8'h00;
im[3208]= 8'h13;
im[3209]= 8'h05;
im[3210]= 8'h85;
im[3211]= 8'h7B;
im[3212]= 8'h33;
im[3213]= 8'h05;
im[3214]= 8'h85;
im[3215]= 8'h00;
im[3216]= 8'h13;
im[3217]= 8'h05;
im[3218]= 8'h05;
im[3219]= 8'h7B;
im[3220]= 8'h33;
im[3221]= 8'h05;
im[3222]= 8'h85;
im[3223]= 8'h00;
im[3224]= 8'h13;
im[3225]= 8'h05;
im[3226]= 8'h85;
im[3227]= 8'h7B;
im[3228]= 8'h33;
im[3229]= 8'h05;
im[3230]= 8'h85;
im[3231]= 8'h00;
im[3232]= 8'h13;
im[3233]= 8'h05;
im[3234]= 8'h05;
im[3235]= 8'h7C;
im[3236]= 8'h33;
im[3237]= 8'h05;
im[3238]= 8'h85;
im[3239]= 8'h00;
im[3240]= 8'h13;
im[3241]= 8'h05;
im[3242]= 8'h85;
im[3243]= 8'h7C;
im[3244]= 8'h33;
im[3245]= 8'h05;
im[3246]= 8'h85;
im[3247]= 8'h00;
im[3248]= 8'h13;
im[3249]= 8'h05;
im[3250]= 8'h04;
im[3251]= 8'h8C;
im[3252]= 8'h13;
im[3253]= 8'h05;
im[3254]= 8'h05;
im[3255]= 8'h7D;
im[3256]= 8'h33;
im[3257]= 8'h05;
im[3258]= 8'h85;
im[3259]= 8'h00;
im[3260]= 8'h83;
im[3261]= 8'h27;
im[3262]= 8'h05;
im[3263]= 8'h00;
im[3264]= 8'h13;
im[3265]= 8'h05;
im[3266]= 8'h45;
im[3267]= 8'h7D;
im[3268]= 8'h33;
im[3269]= 8'h05;
im[3270]= 8'h85;
im[3271]= 8'h00;
im[3272]= 8'h03;
im[3273]= 8'h27;
im[3274]= 8'h05;
im[3275]= 8'h00;
im[3276]= 8'h03;
im[3277]= 8'h25;
im[3278]= 8'h04;
im[3279]= 8'h8C;
im[3280]= 8'h93;
im[3281]= 8'h85;
im[3282]= 8'h45;
im[3283]= 8'h7E;
im[3284]= 8'hB3;
im[3285]= 8'h85;
im[3286]= 8'h85;
im[3287]= 8'h00;
im[3288]= 8'h23;
im[3289]= 8'hA0;
im[3290]= 8'hA5;
im[3291]= 8'h00;
im[3292]= 8'h03;
im[3293]= 8'h25;
im[3294]= 8'h44;
im[3295]= 8'h8C;
im[3296]= 8'h93;
im[3297]= 8'h85;
im[3298]= 8'h05;
im[3299]= 8'h7E;
im[3300]= 8'hB3;
im[3301]= 8'h85;
im[3302]= 8'h85;
im[3303]= 8'h00;
im[3304]= 8'h23;
im[3305]= 8'hA0;
im[3306]= 8'hA5;
im[3307]= 8'h00;
im[3308]= 8'h03;
im[3309]= 8'h25;
im[3310]= 8'h84;
im[3311]= 8'h8C;
im[3312]= 8'h93;
im[3313]= 8'h85;
im[3314]= 8'hC5;
im[3315]= 8'h7D;
im[3316]= 8'hB3;
im[3317]= 8'h85;
im[3318]= 8'h85;
im[3319]= 8'h00;
im[3320]= 8'h23;
im[3321]= 8'hA0;
im[3322]= 8'hA5;
im[3323]= 8'h00;
im[3324]= 8'h03;
im[3325]= 8'h25;
im[3326]= 8'hC4;
im[3327]= 8'h8C;
im[3328]= 8'h93;
im[3329]= 8'h85;
im[3330]= 8'h85;
im[3331]= 8'h7D;
im[3332]= 8'hB3;
im[3333]= 8'h85;
im[3334]= 8'h85;
im[3335]= 8'h00;
im[3336]= 8'h23;
im[3337]= 8'hA0;
im[3338]= 8'hA5;
im[3339]= 8'h00;
im[3340]= 8'h03;
im[3341]= 8'h25;
im[3342]= 8'h04;
im[3343]= 8'hFB;
im[3344]= 8'h83;
im[3345]= 8'h25;
im[3346]= 8'h44;
im[3347]= 8'hFB;
im[3348]= 8'h03;
im[3349]= 8'h26;
im[3350]= 8'h84;
im[3351]= 8'hFB;
im[3352]= 8'h83;
im[3353]= 8'h26;
im[3354]= 8'hC4;
im[3355]= 8'hFB;
im[3356]= 8'h23;
im[3357]= 8'h2E;
im[3358]= 8'hF4;
im[3359]= 8'h88;
im[3360]= 8'h23;
im[3361]= 8'h2C;
im[3362]= 8'hE4;
im[3363]= 8'h88;
im[3364]= 8'h23;
im[3365]= 8'h2A;
im[3366]= 8'hE4;
im[3367]= 8'h88;
im[3368]= 8'h23;
im[3369]= 8'h28;
im[3370]= 8'hE4;
im[3371]= 8'h88;
im[3372]= 8'h23;
im[3373]= 8'h26;
im[3374]= 8'hD4;
im[3375]= 8'h8A;
im[3376]= 8'h23;
im[3377]= 8'h24;
im[3378]= 8'hC4;
im[3379]= 8'h8A;
im[3380]= 8'h23;
im[3381]= 8'h22;
im[3382]= 8'hB4;
im[3383]= 8'h8A;
im[3384]= 8'h23;
im[3385]= 8'h20;
im[3386]= 8'hA4;
im[3387]= 8'h8A;
im[3388]= 8'h13;
im[3389]= 8'h05;
im[3390]= 8'h04;
im[3391]= 8'h8B;
im[3392]= 8'h93;
im[3393]= 8'h05;
im[3394]= 8'h04;
im[3395]= 8'h8A;
im[3396]= 8'h13;
im[3397]= 8'h06;
im[3398]= 8'h04;
im[3399]= 8'h89;
im[3400]= 8'h13;
im[3401]= 8'h05;
im[3402]= 8'h85;
im[3403]= 8'h7D;
im[3404]= 8'h33;
im[3405]= 8'h05;
im[3406]= 8'h85;
im[3407]= 8'h00;
im[3408]= 8'h83;
im[3409]= 8'h28;
im[3410]= 8'h05;
im[3411]= 8'h00;
im[3412]= 8'h13;
im[3413]= 8'h05;
im[3414]= 8'hC5;
im[3415]= 8'h7D;
im[3416]= 8'h33;
im[3417]= 8'h05;
im[3418]= 8'h85;
im[3419]= 8'h00;
im[3420]= 8'h03;
im[3421]= 8'h28;
im[3422]= 8'h05;
im[3423]= 8'h00;
im[3424]= 8'h13;
im[3425]= 8'h05;
im[3426]= 8'h05;
im[3427]= 8'h7E;
im[3428]= 8'h33;
im[3429]= 8'h05;
im[3430]= 8'h85;
im[3431]= 8'h00;
im[3432]= 8'h83;
im[3433]= 8'h27;
im[3434]= 8'h05;
im[3435]= 8'h00;
im[3436]= 8'h13;
im[3437]= 8'h05;
im[3438]= 8'h45;
im[3439]= 8'h7E;
im[3440]= 8'h33;
im[3441]= 8'h05;
im[3442]= 8'h85;
im[3443]= 8'h00;
im[3444]= 8'h03;
im[3445]= 8'h27;
im[3446]= 8'h05;
im[3447]= 8'h00;
im[3448]= 8'h03;
im[3449]= 8'h25;
im[3450]= 8'h04;
im[3451]= 8'h8B;
im[3452]= 8'h83;
im[3453]= 8'h25;
im[3454]= 8'h44;
im[3455]= 8'h8B;
im[3456]= 8'h03;
im[3457]= 8'h26;
im[3458]= 8'h84;
im[3459]= 8'h8B;
im[3460]= 8'h83;
im[3461]= 8'h26;
im[3462]= 8'hC4;
im[3463]= 8'h8B;
im[3464]= 8'h23;
im[3465]= 8'h2E;
im[3466]= 8'h14;
im[3467]= 8'h87;
im[3468]= 8'h23;
im[3469]= 8'h2C;
im[3470]= 8'h04;
im[3471]= 8'h87;
im[3472]= 8'h23;
im[3473]= 8'h2A;
im[3474]= 8'hF4;
im[3475]= 8'h86;
im[3476]= 8'h23;
im[3477]= 8'h28;
im[3478]= 8'hE4;
im[3479]= 8'h86;
im[3480]= 8'h23;
im[3481]= 8'h26;
im[3482]= 8'hD4;
im[3483]= 8'h86;
im[3484]= 8'h23;
im[3485]= 8'h24;
im[3486]= 8'hC4;
im[3487]= 8'h86;
im[3488]= 8'h23;
im[3489]= 8'h22;
im[3490]= 8'hB4;
im[3491]= 8'h86;
im[3492]= 8'h23;
im[3493]= 8'h20;
im[3494]= 8'hA4;
im[3495]= 8'h86;
im[3496]= 8'h13;
im[3497]= 8'h05;
im[3498]= 8'h04;
im[3499]= 8'h88;
im[3500]= 8'h93;
im[3501]= 8'h05;
im[3502]= 8'h04;
im[3503]= 8'h87;
im[3504]= 8'h13;
im[3505]= 8'h06;
im[3506]= 8'h04;
im[3507]= 8'h86;
im[3508]= 8'h03;
im[3509]= 8'h25;
im[3510]= 8'h04;
im[3511]= 8'h88;
im[3512]= 8'h83;
im[3513]= 8'h25;
im[3514]= 8'h44;
im[3515]= 8'h88;
im[3516]= 8'h03;
im[3517]= 8'h26;
im[3518]= 8'h84;
im[3519]= 8'h88;
im[3520]= 8'h83;
im[3521]= 8'h26;
im[3522]= 8'hC4;
im[3523]= 8'h88;
im[3524]= 8'h23;
im[3525]= 8'h2E;
im[3526]= 8'hD4;
im[3527]= 8'h84;
im[3528]= 8'h23;
im[3529]= 8'h2C;
im[3530]= 8'hC4;
im[3531]= 8'h84;
im[3532]= 8'h23;
im[3533]= 8'h2A;
im[3534]= 8'hB4;
im[3535]= 8'h84;
im[3536]= 8'h23;
im[3537]= 8'h28;
im[3538]= 8'hA4;
im[3539]= 8'h84;
im[3540]= 8'h13;
im[3541]= 8'h05;
im[3542]= 8'h04;
im[3543]= 8'h85;
im[3544]= 8'h03;
im[3545]= 8'h25;
im[3546]= 8'h84;
im[3547]= 8'hFC;
im[3548]= 8'h6F;
im[3549]= 8'h00;
im[3550]= 8'h00;
im[3551]= 8'h3C;
im[3552]= 8'h83;
im[3553]= 8'h25;
im[3554]= 8'hC4;
im[3555]= 8'hFC;
im[3556]= 8'h13;
im[3557]= 8'h05;
im[3558]= 8'h10;
im[3559]= 8'h00;
im[3560]= 8'h13;
im[3561]= 8'h06;
im[3562]= 8'h86;
im[3563]= 8'h73;
im[3564]= 8'h33;
im[3565]= 8'h06;
im[3566]= 8'h86;
im[3567]= 8'h00;
im[3568]= 8'h23;
im[3569]= 8'h20;
im[3570]= 8'hA6;
im[3571]= 8'h00;
im[3572]= 8'h23;
im[3573]= 8'hA0;
im[3574]= 8'hA5;
im[3575]= 8'h00;
im[3576]= 8'h13;
im[3577]= 8'h05;
im[3578]= 8'h85;
im[3579]= 8'h70;
im[3580]= 8'h33;
im[3581]= 8'h05;
im[3582]= 8'h85;
im[3583]= 8'h00;
im[3584]= 8'h03;
im[3585]= 8'h25;
im[3586]= 8'h04;
im[3587]= 8'hF7;
im[3588]= 8'h83;
im[3589]= 8'h25;
im[3590]= 8'h44;
im[3591]= 8'hF7;
im[3592]= 8'h03;
im[3593]= 8'h26;
im[3594]= 8'h84;
im[3595]= 8'hF7;
im[3596]= 8'h83;
im[3597]= 8'h26;
im[3598]= 8'hC4;
im[3599]= 8'hF7;
im[3600]= 8'h23;
im[3601]= 8'h26;
im[3602]= 8'hD4;
im[3603]= 8'hBE;
im[3604]= 8'h23;
im[3605]= 8'h24;
im[3606]= 8'hC4;
im[3607]= 8'hBE;
im[3608]= 8'h23;
im[3609]= 8'h22;
im[3610]= 8'hB4;
im[3611]= 8'hBE;
im[3612]= 8'h23;
im[3613]= 8'h20;
im[3614]= 8'hA4;
im[3615]= 8'hBE;
im[3616]= 8'h13;
im[3617]= 8'h05;
im[3618]= 8'h04;
im[3619]= 8'hBE;
im[3620]= 8'h13;
im[3621]= 8'h05;
im[3622]= 8'h85;
im[3623]= 8'h70;
im[3624]= 8'h33;
im[3625]= 8'h05;
im[3626]= 8'h85;
im[3627]= 8'h00;
im[3628]= 8'h03;
im[3629]= 8'h25;
im[3630]= 8'h84;
im[3631]= 8'hFC;
im[3632]= 8'h03;
im[3633]= 8'h25;
im[3634]= 8'h04;
im[3635]= 8'hF8;
im[3636]= 8'h93;
im[3637]= 8'h85;
im[3638]= 8'h05;
im[3639]= 8'h72;
im[3640]= 8'hB3;
im[3641]= 8'h85;
im[3642]= 8'h85;
im[3643]= 8'h00;
im[3644]= 8'h23;
im[3645]= 8'hA0;
im[3646]= 8'hA5;
im[3647]= 8'h00;
im[3648]= 8'h03;
im[3649]= 8'h25;
im[3650]= 8'h44;
im[3651]= 8'hF8;
im[3652]= 8'h93;
im[3653]= 8'h85;
im[3654]= 8'hC5;
im[3655]= 8'h71;
im[3656]= 8'hB3;
im[3657]= 8'h85;
im[3658]= 8'h85;
im[3659]= 8'h00;
im[3660]= 8'h23;
im[3661]= 8'hA0;
im[3662]= 8'hA5;
im[3663]= 8'h00;
im[3664]= 8'h03;
im[3665]= 8'h25;
im[3666]= 8'h84;
im[3667]= 8'hF8;
im[3668]= 8'h93;
im[3669]= 8'h85;
im[3670]= 8'h85;
im[3671]= 8'h71;
im[3672]= 8'hB3;
im[3673]= 8'h85;
im[3674]= 8'h85;
im[3675]= 8'h00;
im[3676]= 8'h23;
im[3677]= 8'hA0;
im[3678]= 8'hA5;
im[3679]= 8'h00;
im[3680]= 8'h03;
im[3681]= 8'h25;
im[3682]= 8'hC4;
im[3683]= 8'hF8;
im[3684]= 8'h93;
im[3685]= 8'h85;
im[3686]= 8'h45;
im[3687]= 8'h71;
im[3688]= 8'hB3;
im[3689]= 8'h85;
im[3690]= 8'h85;
im[3691]= 8'h00;
im[3692]= 8'h23;
im[3693]= 8'hA0;
im[3694]= 8'hA5;
im[3695]= 8'h00;
im[3696]= 8'h03;
im[3697]= 8'h25;
im[3698]= 8'h84;
im[3699]= 8'hFC;
im[3700]= 8'h93;
im[3701]= 8'h85;
im[3702]= 8'h45;
im[3703]= 8'h73;
im[3704]= 8'hB3;
im[3705]= 8'h85;
im[3706]= 8'h85;
im[3707]= 8'h00;
im[3708]= 8'h23;
im[3709]= 8'hA0;
im[3710]= 8'hA5;
im[3711]= 8'h00;
im[3712]= 8'h13;
im[3713]= 8'h05;
im[3714]= 8'h04;
im[3715]= 8'hB6;
im[3716]= 8'h13;
im[3717]= 8'h05;
im[3718]= 8'h45;
im[3719]= 8'h71;
im[3720]= 8'h33;
im[3721]= 8'h05;
im[3722]= 8'h85;
im[3723]= 8'h00;
im[3724]= 8'h83;
im[3725]= 8'h28;
im[3726]= 8'h05;
im[3727]= 8'h00;
im[3728]= 8'h13;
im[3729]= 8'h05;
im[3730]= 8'h85;
im[3731]= 8'h71;
im[3732]= 8'h33;
im[3733]= 8'h05;
im[3734]= 8'h85;
im[3735]= 8'h00;
im[3736]= 8'h03;
im[3737]= 8'h28;
im[3738]= 8'h05;
im[3739]= 8'h00;
im[3740]= 8'h13;
im[3741]= 8'h05;
im[3742]= 8'hC5;
im[3743]= 8'h71;
im[3744]= 8'h33;
im[3745]= 8'h05;
im[3746]= 8'h85;
im[3747]= 8'h00;
im[3748]= 8'h83;
im[3749]= 8'h27;
im[3750]= 8'h05;
im[3751]= 8'h00;
im[3752]= 8'h13;
im[3753]= 8'h05;
im[3754]= 8'h05;
im[3755]= 8'h72;
im[3756]= 8'h33;
im[3757]= 8'h05;
im[3758]= 8'h85;
im[3759]= 8'h00;
im[3760]= 8'h03;
im[3761]= 8'h27;
im[3762]= 8'h05;
im[3763]= 8'h00;
im[3764]= 8'h03;
im[3765]= 8'h25;
im[3766]= 8'h04;
im[3767]= 8'hB6;
im[3768]= 8'h93;
im[3769]= 8'h85;
im[3770]= 8'h05;
im[3771]= 8'h73;
im[3772]= 8'hB3;
im[3773]= 8'h85;
im[3774]= 8'h85;
im[3775]= 8'h00;
im[3776]= 8'h23;
im[3777]= 8'hA0;
im[3778]= 8'hA5;
im[3779]= 8'h00;
im[3780]= 8'h83;
im[3781]= 8'h25;
im[3782]= 8'h44;
im[3783]= 8'hB6;
im[3784]= 8'h13;
im[3785]= 8'h06;
im[3786]= 8'hC6;
im[3787]= 8'h72;
im[3788]= 8'h33;
im[3789]= 8'h06;
im[3790]= 8'h86;
im[3791]= 8'h00;
im[3792]= 8'h23;
im[3793]= 8'h20;
im[3794]= 8'hB6;
im[3795]= 8'h00;
im[3796]= 8'h03;
im[3797]= 8'h26;
im[3798]= 8'h84;
im[3799]= 8'hB6;
im[3800]= 8'h93;
im[3801]= 8'h86;
im[3802]= 8'h86;
im[3803]= 8'h72;
im[3804]= 8'hB3;
im[3805]= 8'h86;
im[3806]= 8'h86;
im[3807]= 8'h00;
im[3808]= 8'h23;
im[3809]= 8'hA0;
im[3810]= 8'hC6;
im[3811]= 8'h00;
im[3812]= 8'h83;
im[3813]= 8'h26;
im[3814]= 8'hC4;
im[3815]= 8'hB6;
im[3816]= 8'h93;
im[3817]= 8'h82;
im[3818]= 8'h42;
im[3819]= 8'h72;
im[3820]= 8'hB3;
im[3821]= 8'h82;
im[3822]= 8'h82;
im[3823]= 8'h00;
im[3824]= 8'h23;
im[3825]= 8'hA0;
im[3826]= 8'hD2;
im[3827]= 8'h00;
im[3828]= 8'h23;
im[3829]= 8'h26;
im[3830]= 8'h14;
im[3831]= 8'hBD;
im[3832]= 8'h23;
im[3833]= 8'h24;
im[3834]= 8'h04;
im[3835]= 8'hBD;
im[3836]= 8'h23;
im[3837]= 8'h22;
im[3838]= 8'hF4;
im[3839]= 8'hBC;
im[3840]= 8'h23;
im[3841]= 8'h20;
im[3842]= 8'hE4;
im[3843]= 8'hBC;
im[3844]= 8'h23;
im[3845]= 8'h2E;
im[3846]= 8'hD4;
im[3847]= 8'hBA;
im[3848]= 8'h23;
im[3849]= 8'h2C;
im[3850]= 8'hC4;
im[3851]= 8'hBA;
im[3852]= 8'h23;
im[3853]= 8'h2A;
im[3854]= 8'hB4;
im[3855]= 8'hBA;
im[3856]= 8'h23;
im[3857]= 8'h28;
im[3858]= 8'hA4;
im[3859]= 8'hBA;
im[3860]= 8'h13;
im[3861]= 8'h05;
im[3862]= 8'h04;
im[3863]= 8'hBD;
im[3864]= 8'h93;
im[3865]= 8'h05;
im[3866]= 8'h04;
im[3867]= 8'hBC;
im[3868]= 8'h13;
im[3869]= 8'h06;
im[3870]= 8'h04;
im[3871]= 8'hBB;
im[3872]= 8'h13;
im[3873]= 8'h05;
im[3874]= 8'h45;
im[3875]= 8'h72;
im[3876]= 8'h33;
im[3877]= 8'h05;
im[3878]= 8'h85;
im[3879]= 8'h00;
im[3880]= 8'h83;
im[3881]= 8'h28;
im[3882]= 8'h05;
im[3883]= 8'h00;
im[3884]= 8'h13;
im[3885]= 8'h05;
im[3886]= 8'h85;
im[3887]= 8'h72;
im[3888]= 8'h33;
im[3889]= 8'h05;
im[3890]= 8'h85;
im[3891]= 8'h00;
im[3892]= 8'h03;
im[3893]= 8'h28;
im[3894]= 8'h05;
im[3895]= 8'h00;
im[3896]= 8'h13;
im[3897]= 8'h05;
im[3898]= 8'hC5;
im[3899]= 8'h72;
im[3900]= 8'h33;
im[3901]= 8'h05;
im[3902]= 8'h85;
im[3903]= 8'h00;
im[3904]= 8'h83;
im[3905]= 8'h27;
im[3906]= 8'h05;
im[3907]= 8'h00;
im[3908]= 8'h13;
im[3909]= 8'h05;
im[3910]= 8'h05;
im[3911]= 8'h73;
im[3912]= 8'h33;
im[3913]= 8'h05;
im[3914]= 8'h85;
im[3915]= 8'h00;
im[3916]= 8'h03;
im[3917]= 8'h27;
im[3918]= 8'h05;
im[3919]= 8'h00;
im[3920]= 8'h03;
im[3921]= 8'h25;
im[3922]= 8'h04;
im[3923]= 8'hBD;
im[3924]= 8'h83;
im[3925]= 8'h25;
im[3926]= 8'h44;
im[3927]= 8'hBD;
im[3928]= 8'h03;
im[3929]= 8'h26;
im[3930]= 8'h84;
im[3931]= 8'hBD;
im[3932]= 8'h83;
im[3933]= 8'h26;
im[3934]= 8'hC4;
im[3935]= 8'hBD;
im[3936]= 8'h23;
im[3937]= 8'h2E;
im[3938]= 8'h14;
im[3939]= 8'hB9;
im[3940]= 8'h23;
im[3941]= 8'h2C;
im[3942]= 8'h04;
im[3943]= 8'hB9;
im[3944]= 8'h23;
im[3945]= 8'h2A;
im[3946]= 8'hF4;
im[3947]= 8'hB8;
im[3948]= 8'h23;
im[3949]= 8'h28;
im[3950]= 8'hE4;
im[3951]= 8'hB8;
im[3952]= 8'h23;
im[3953]= 8'h26;
im[3954]= 8'hD4;
im[3955]= 8'hB8;
im[3956]= 8'h23;
im[3957]= 8'h24;
im[3958]= 8'hC4;
im[3959]= 8'hB8;
im[3960]= 8'h23;
im[3961]= 8'h22;
im[3962]= 8'hB4;
im[3963]= 8'hB8;
im[3964]= 8'h23;
im[3965]= 8'h20;
im[3966]= 8'hA4;
im[3967]= 8'hB8;
im[3968]= 8'h13;
im[3969]= 8'h05;
im[3970]= 8'h04;
im[3971]= 8'hBA;
im[3972]= 8'h93;
im[3973]= 8'h05;
im[3974]= 8'h04;
im[3975]= 8'hB9;
im[3976]= 8'h13;
im[3977]= 8'h06;
im[3978]= 8'h04;
im[3979]= 8'hB8;
im[3980]= 8'h03;
im[3981]= 8'h25;
im[3982]= 8'h04;
im[3983]= 8'hBA;
im[3984]= 8'h83;
im[3985]= 8'h25;
im[3986]= 8'h44;
im[3987]= 8'hBA;
im[3988]= 8'h03;
im[3989]= 8'h26;
im[3990]= 8'h84;
im[3991]= 8'hBA;
im[3992]= 8'h83;
im[3993]= 8'h26;
im[3994]= 8'hC4;
im[3995]= 8'hBA;
im[3996]= 8'h23;
im[3997]= 8'h2E;
im[3998]= 8'hD4;
im[3999]= 8'hB6;
im[4000]= 8'h23;
im[4001]= 8'h2C;
im[4002]= 8'hC4;
im[4003]= 8'hB6;
im[4004]= 8'h23;
im[4005]= 8'h2A;
im[4006]= 8'hB4;
im[4007]= 8'hB6;
im[4008]= 8'h23;
im[4009]= 8'h28;
im[4010]= 8'hA4;
im[4011]= 8'hB6;
im[4012]= 8'h13;
im[4013]= 8'h05;
im[4014]= 8'h04;
im[4015]= 8'hB7;
im[4016]= 8'h13;
im[4017]= 8'h05;
im[4018]= 8'h45;
im[4019]= 8'h73;
im[4020]= 8'h33;
im[4021]= 8'h05;
im[4022]= 8'h85;
im[4023]= 8'h00;
im[4024]= 8'h03;
im[4025]= 8'h25;
im[4026]= 8'h05;
im[4027]= 8'h00;
im[4028]= 8'h03;
im[4029]= 8'h25;
im[4030]= 8'h04;
im[4031]= 8'hF7;
im[4032]= 8'h83;
im[4033]= 8'h25;
im[4034]= 8'h44;
im[4035]= 8'hF7;
im[4036]= 8'h03;
im[4037]= 8'h26;
im[4038]= 8'h84;
im[4039]= 8'hF7;
im[4040]= 8'h83;
im[4041]= 8'h26;
im[4042]= 8'hC4;
im[4043]= 8'hF7;
im[4044]= 8'h93;
im[4045]= 8'h87;
im[4046]= 8'hC7;
im[4047]= 8'h73;
im[4048]= 8'hB3;
im[4049]= 8'h87;
im[4050]= 8'h87;
im[4051]= 8'h00;
im[4052]= 8'h23;
im[4053]= 8'hA0;
im[4054]= 8'hE7;
im[4055]= 8'h00;
im[4056]= 8'h23;
im[4057]= 8'h26;
im[4058]= 8'hE4;
im[4059]= 8'hB4;
im[4060]= 8'h23;
im[4061]= 8'h24;
im[4062]= 8'hE4;
im[4063]= 8'hB4;
im[4064]= 8'h23;
im[4065]= 8'h22;
im[4066]= 8'hE4;
im[4067]= 8'hB4;
im[4068]= 8'h23;
im[4069]= 8'h20;
im[4070]= 8'hE4;
im[4071]= 8'hB4;
im[4072]= 8'h23;
im[4073]= 8'h2E;
im[4074]= 8'hD4;
im[4075]= 8'hB4;
im[4076]= 8'h23;
im[4077]= 8'h2C;
im[4078]= 8'hC4;
im[4079]= 8'hB4;
im[4080]= 8'h23;
im[4081]= 8'h2A;
im[4082]= 8'hB4;
im[4083]= 8'hB4;
im[4084]= 8'h23;
im[4085]= 8'h28;
im[4086]= 8'hA4;
im[4087]= 8'hB4;
im[4088]= 8'h13;
im[4089]= 8'h05;
im[4090]= 8'h04;
im[4091]= 8'hB5;
im[4092]= 8'h93;
im[4093]= 8'h05;
im[4094]= 8'h04;
im[4095]= 8'hB4;
im[4096]= 8'h93;
im[4097]= 8'h85;
im[4098]= 8'h85;
im[4099]= 8'h73;
im[4100]= 8'hB3;
im[4101]= 8'h85;
im[4102]= 8'h85;
im[4103]= 8'h00;
im[4104]= 8'h03;
im[4105]= 8'hA6;
im[4106]= 8'h05;
im[4107]= 8'h00;
im[4108]= 8'h93;
im[4109]= 8'h85;
im[4110]= 8'hC5;
im[4111]= 8'h73;
im[4112]= 8'hB3;
im[4113]= 8'h85;
im[4114]= 8'h85;
im[4115]= 8'h00;
im[4116]= 8'h83;
im[4117]= 8'hA5;
im[4118]= 8'h05;
im[4119]= 8'h00;
im[4120]= 8'h93;
im[4121]= 8'h06;
im[4122]= 8'hF0;
im[4123]= 8'hFF;
im[4124]= 8'h13;
im[4125]= 8'h07;
im[4126]= 8'h07;
im[4127]= 8'h74;
im[4128]= 8'h33;
im[4129]= 8'h07;
im[4130]= 8'h87;
im[4131]= 8'h00;
im[4132]= 8'h23;
im[4133]= 8'h20;
im[4134]= 8'hD7;
im[4135]= 8'h00;
im[4136]= 8'h93;
im[4137]= 8'h86;
im[4138]= 8'h46;
im[4139]= 8'h74;
im[4140]= 8'hB3;
im[4141]= 8'h86;
im[4142]= 8'h86;
im[4143]= 8'h00;
im[4144]= 8'h23;
im[4145]= 8'hA0;
im[4146]= 8'hC6;
im[4147]= 8'h00;
im[4148]= 8'h63;
im[4149]= 8'h4E;
im[4150]= 8'hB5;
im[4151]= 8'h00;
im[4152]= 8'h13;
im[4153]= 8'h05;
im[4154]= 8'h05;
im[4155]= 8'h74;
im[4156]= 8'h33;
im[4157]= 8'h05;
im[4158]= 8'h85;
im[4159]= 8'h00;
im[4160]= 8'h03;
im[4161]= 8'h25;
im[4162]= 8'h05;
im[4163]= 8'h00;
im[4164]= 8'h93;
im[4165]= 8'h85;
im[4166]= 8'h45;
im[4167]= 8'h74;
im[4168]= 8'hB3;
im[4169]= 8'h85;
im[4170]= 8'h85;
im[4171]= 8'h00;
im[4172]= 8'h23;
im[4173]= 8'hA0;
im[4174]= 8'hA5;
im[4175]= 8'h00;
im[4176]= 8'h13;
im[4177]= 8'h05;
im[4178]= 8'hC5;
im[4179]= 8'h73;
im[4180]= 8'h33;
im[4181]= 8'h05;
im[4182]= 8'h85;
im[4183]= 8'h00;
im[4184]= 8'h03;
im[4185]= 8'h27;
im[4186]= 8'h05;
im[4187]= 8'h00;
im[4188]= 8'h13;
im[4189]= 8'h05;
im[4190]= 8'h45;
im[4191]= 8'h74;
im[4192]= 8'h33;
im[4193]= 8'h05;
im[4194]= 8'h85;
im[4195]= 8'h00;
im[4196]= 8'h03;
im[4197]= 8'h25;
im[4198]= 8'h05;
im[4199]= 8'h00;
im[4200]= 8'h03;
im[4201]= 8'h25;
im[4202]= 8'h84;
im[4203]= 8'hFC;
im[4204]= 8'h03;
im[4205]= 8'h25;
im[4206]= 8'h04;
im[4207]= 8'hFB;
im[4208]= 8'h83;
im[4209]= 8'h25;
im[4210]= 8'h44;
im[4211]= 8'hFB;
im[4212]= 8'h03;
im[4213]= 8'h26;
im[4214]= 8'h84;
im[4215]= 8'hFB;
im[4216]= 8'h83;
im[4217]= 8'h26;
im[4218]= 8'hC4;
im[4219]= 8'hFB;
im[4220]= 8'h23;
im[4221]= 8'h2E;
im[4222]= 8'hF4;
im[4223]= 8'hB0;
im[4224]= 8'h23;
im[4225]= 8'h2C;
im[4226]= 8'hE4;
im[4227]= 8'hB0;
im[4228]= 8'h23;
im[4229]= 8'h2A;
im[4230]= 8'hE4;
im[4231]= 8'hB0;
im[4232]= 8'h23;
im[4233]= 8'h28;
im[4234]= 8'hE4;
im[4235]= 8'hB0;
im[4236]= 8'h23;
im[4237]= 8'h26;
im[4238]= 8'hD4;
im[4239]= 8'hB2;
im[4240]= 8'h23;
im[4241]= 8'h24;
im[4242]= 8'hC4;
im[4243]= 8'hB2;
im[4244]= 8'h23;
im[4245]= 8'h22;
im[4246]= 8'hB4;
im[4247]= 8'hB2;
im[4248]= 8'h23;
im[4249]= 8'h20;
im[4250]= 8'hA4;
im[4251]= 8'hB2;
im[4252]= 8'h13;
im[4253]= 8'h05;
im[4254]= 8'h04;
im[4255]= 8'hB3;
im[4256]= 8'h93;
im[4257]= 8'h05;
im[4258]= 8'h04;
im[4259]= 8'hB2;
im[4260]= 8'h13;
im[4261]= 8'h06;
im[4262]= 8'h04;
im[4263]= 8'hB1;
im[4264]= 8'h03;
im[4265]= 8'h25;
im[4266]= 8'h04;
im[4267]= 8'hB3;
im[4268]= 8'h93;
im[4269]= 8'h85;
im[4270]= 8'h05;
im[4271]= 8'h70;
im[4272]= 8'hB3;
im[4273]= 8'h85;
im[4274]= 8'h85;
im[4275]= 8'h00;
im[4276]= 8'h23;
im[4277]= 8'hA0;
im[4278]= 8'hA5;
im[4279]= 8'h00;
im[4280]= 8'h03;
im[4281]= 8'h25;
im[4282]= 8'h44;
im[4283]= 8'hB3;
im[4284]= 8'h93;
im[4285]= 8'h85;
im[4286]= 8'hC5;
im[4287]= 8'h6F;
im[4288]= 8'hB3;
im[4289]= 8'h85;
im[4290]= 8'h85;
im[4291]= 8'h00;
im[4292]= 8'h23;
im[4293]= 8'hA0;
im[4294]= 8'hA5;
im[4295]= 8'h00;
im[4296]= 8'h03;
im[4297]= 8'h25;
im[4298]= 8'h84;
im[4299]= 8'hB3;
im[4300]= 8'h93;
im[4301]= 8'h85;
im[4302]= 8'h85;
im[4303]= 8'h6F;
im[4304]= 8'hB3;
im[4305]= 8'h85;
im[4306]= 8'h85;
im[4307]= 8'h00;
im[4308]= 8'h23;
im[4309]= 8'hA0;
im[4310]= 8'hA5;
im[4311]= 8'h00;
im[4312]= 8'h03;
im[4313]= 8'h25;
im[4314]= 8'hC4;
im[4315]= 8'hB3;
im[4316]= 8'h93;
im[4317]= 8'h85;
im[4318]= 8'h45;
im[4319]= 8'h6F;
im[4320]= 8'hB3;
im[4321]= 8'h85;
im[4322]= 8'h85;
im[4323]= 8'h00;
im[4324]= 8'h23;
im[4325]= 8'hA0;
im[4326]= 8'hA5;
im[4327]= 8'h00;
im[4328]= 8'h03;
im[4329]= 8'h25;
im[4330]= 8'h84;
im[4331]= 8'hFC;
im[4332]= 8'h93;
im[4333]= 8'h85;
im[4334]= 8'h45;
im[4335]= 8'h70;
im[4336]= 8'hB3;
im[4337]= 8'h85;
im[4338]= 8'h85;
im[4339]= 8'h00;
im[4340]= 8'h23;
im[4341]= 8'hA0;
im[4342]= 8'hA5;
im[4343]= 8'h00;
im[4344]= 8'h13;
im[4345]= 8'h05;
im[4346]= 8'h04;
im[4347]= 8'hAC;
im[4348]= 8'h13;
im[4349]= 8'h05;
im[4350]= 8'h45;
im[4351]= 8'h6F;
im[4352]= 8'h33;
im[4353]= 8'h05;
im[4354]= 8'h85;
im[4355]= 8'h00;
im[4356]= 8'h83;
im[4357]= 8'h28;
im[4358]= 8'h05;
im[4359]= 8'h00;
im[4360]= 8'h13;
im[4361]= 8'h05;
im[4362]= 8'h85;
im[4363]= 8'h6F;
im[4364]= 8'h33;
im[4365]= 8'h05;
im[4366]= 8'h85;
im[4367]= 8'h00;
im[4368]= 8'h03;
im[4369]= 8'h28;
im[4370]= 8'h05;
im[4371]= 8'h00;
im[4372]= 8'h13;
im[4373]= 8'h05;
im[4374]= 8'hC5;
im[4375]= 8'h6F;
im[4376]= 8'h33;
im[4377]= 8'h05;
im[4378]= 8'h85;
im[4379]= 8'h00;
im[4380]= 8'h83;
im[4381]= 8'h27;
im[4382]= 8'h05;
im[4383]= 8'h00;
im[4384]= 8'h13;
im[4385]= 8'h05;
im[4386]= 8'h05;
im[4387]= 8'h70;
im[4388]= 8'h33;
im[4389]= 8'h05;
im[4390]= 8'h85;
im[4391]= 8'h00;
im[4392]= 8'h03;
im[4393]= 8'h27;
im[4394]= 8'h05;
im[4395]= 8'h00;
im[4396]= 8'h03;
im[4397]= 8'h25;
im[4398]= 8'h04;
im[4399]= 8'hAC;
im[4400]= 8'h83;
im[4401]= 8'h25;
im[4402]= 8'h44;
im[4403]= 8'hAC;
im[4404]= 8'h03;
im[4405]= 8'h26;
im[4406]= 8'h84;
im[4407]= 8'hAC;
im[4408]= 8'h83;
im[4409]= 8'h26;
im[4410]= 8'hC4;
im[4411]= 8'hAC;
im[4412]= 8'h23;
im[4413]= 8'h26;
im[4414]= 8'h14;
im[4415]= 8'hAF;
im[4416]= 8'h23;
im[4417]= 8'h24;
im[4418]= 8'h04;
im[4419]= 8'hAF;
im[4420]= 8'h23;
im[4421]= 8'h22;
im[4422]= 8'hF4;
im[4423]= 8'hAE;
im[4424]= 8'h23;
im[4425]= 8'h20;
im[4426]= 8'hE4;
im[4427]= 8'hAE;
im[4428]= 8'h23;
im[4429]= 8'h2E;
im[4430]= 8'hD4;
im[4431]= 8'hAE;
im[4432]= 8'h23;
im[4433]= 8'h2C;
im[4434]= 8'hC4;
im[4435]= 8'hAE;
im[4436]= 8'h23;
im[4437]= 8'h2A;
im[4438]= 8'hB4;
im[4439]= 8'hAE;
im[4440]= 8'h23;
im[4441]= 8'h28;
im[4442]= 8'hA4;
im[4443]= 8'hAE;
im[4444]= 8'h13;
im[4445]= 8'h05;
im[4446]= 8'h04;
im[4447]= 8'hB0;
im[4448]= 8'h93;
im[4449]= 8'h05;
im[4450]= 8'h04;
im[4451]= 8'hAF;
im[4452]= 8'h13;
im[4453]= 8'h06;
im[4454]= 8'h04;
im[4455]= 8'hAE;
im[4456]= 8'h03;
im[4457]= 8'h25;
im[4458]= 8'h04;
im[4459]= 8'hB0;
im[4460]= 8'h83;
im[4461]= 8'h25;
im[4462]= 8'h44;
im[4463]= 8'hB0;
im[4464]= 8'h03;
im[4465]= 8'h26;
im[4466]= 8'h84;
im[4467]= 8'hB0;
im[4468]= 8'h83;
im[4469]= 8'h26;
im[4470]= 8'hC4;
im[4471]= 8'hB0;
im[4472]= 8'h23;
im[4473]= 8'h2E;
im[4474]= 8'hD4;
im[4475]= 8'hAC;
im[4476]= 8'h23;
im[4477]= 8'h2C;
im[4478]= 8'hC4;
im[4479]= 8'hAC;
im[4480]= 8'h23;
im[4481]= 8'h2A;
im[4482]= 8'hB4;
im[4483]= 8'hAC;
im[4484]= 8'h23;
im[4485]= 8'h28;
im[4486]= 8'hA4;
im[4487]= 8'hAC;
im[4488]= 8'h13;
im[4489]= 8'h05;
im[4490]= 8'h04;
im[4491]= 8'hAD;
im[4492]= 8'h13;
im[4493]= 8'h05;
im[4494]= 8'h45;
im[4495]= 8'h70;
im[4496]= 8'h33;
im[4497]= 8'h05;
im[4498]= 8'h85;
im[4499]= 8'h00;
im[4500]= 8'h03;
im[4501]= 8'h25;
im[4502]= 8'h05;
im[4503]= 8'h00;
im[4504]= 8'h6F;
im[4505]= 8'h00;
im[4506]= 8'h40;
im[4507]= 8'h00;
im[4508]= 8'h13;
im[4509]= 8'h01;
im[4510]= 8'h01;
im[4511]= 8'h12;
im[4512]= 8'h03;
im[4513]= 8'h24;
im[4514]= 8'h81;
im[4515]= 8'h7E;
im[4516]= 8'h83;
im[4517]= 8'h20;
im[4518]= 8'hC1;
im[4519]= 8'h7E;
im[4520]= 8'h13;
im[4521]= 8'h01;
im[4522]= 8'h01;
im[4523]= 8'h7F;
im[4524]= 8'h13;
im[4525]= 8'h01;
im[4526]= 8'h01;
im[4527]= 8'hF4;
im[4528]= 8'h23;
im[4529]= 8'h2E;
im[4530]= 8'h11;
im[4531]= 8'h0A;
im[4532]= 8'h23;
im[4533]= 8'h2C;
im[4534]= 8'h81;
im[4535]= 8'h0A;
im[4536]= 8'h13;
im[4537]= 8'h04;
im[4538]= 8'h01;
im[4539]= 8'h0C;
im[4540]= 8'h23;
im[4541]= 8'h22;
im[4542]= 8'hA4;
im[4543]= 8'hF8;
im[4544]= 8'h23;
im[4545]= 8'h2A;
im[4546]= 8'hA4;
im[4547]= 8'hFE;
im[4548]= 8'h23;
im[4549]= 8'h26;
im[4550]= 8'hB4;
im[4551]= 8'hFE;
im[4552]= 8'h23;
im[4553]= 8'h24;
im[4554]= 8'hA4;
im[4555]= 8'hFE;
im[4556]= 8'h23;
im[4557]= 8'h22;
im[4558]= 8'hB4;
im[4559]= 8'hFE;
im[4560]= 8'h23;
im[4561]= 8'h20;
im[4562]= 8'hA4;
im[4563]= 8'hFE;
im[4564]= 8'h23;
im[4565]= 8'h2E;
im[4566]= 8'hB4;
im[4567]= 8'hFC;
im[4568]= 8'h23;
im[4569]= 8'h2C;
im[4570]= 8'hA4;
im[4571]= 8'hFC;
im[4572]= 8'h23;
im[4573]= 8'h2A;
im[4574]= 8'hB4;
im[4575]= 8'hFC;
im[4576]= 8'h23;
im[4577]= 8'h28;
im[4578]= 8'hA4;
im[4579]= 8'hFC;
im[4580]= 8'h93;
im[4581]= 8'h85;
im[4582]= 8'h95;
im[4583]= 8'h16;
im[4584]= 8'h23;
im[4585]= 8'h22;
im[4586]= 8'hB4;
im[4587]= 8'hFA;
im[4588]= 8'h23;
im[4589]= 8'h2A;
im[4590]= 8'hA4;
im[4591]= 8'hF8;
im[4592]= 8'h13;
im[4593]= 8'h05;
im[4594]= 8'hC4;
im[4595]= 8'hFA;
im[4596]= 8'h93;
im[4597]= 8'h05;
im[4598]= 8'h84;
im[4599]= 8'hFB;
im[4600]= 8'h03;
im[4601]= 8'h25;
im[4602]= 8'h44;
im[4603]= 8'hF8;
im[4604]= 8'h23;
im[4605]= 8'h24;
im[4606]= 8'hA4;
im[4607]= 8'hFA;
im[4608]= 8'h6F;
im[4609]= 8'h00;
im[4610]= 8'h40;
im[4611]= 8'h00;
im[4612]= 8'h03;
im[4613]= 8'h25;
im[4614]= 8'h84;
im[4615]= 8'hFA;
im[4616]= 8'h83;
im[4617]= 8'h25;
im[4618]= 8'hC4;
im[4619]= 8'hFA;
im[4620]= 8'h63;
im[4621]= 8'h5A;
im[4622]= 8'hB5;
im[4623]= 8'h02;
im[4624]= 8'h6F;
im[4625]= 8'h00;
im[4626]= 8'h40;
im[4627]= 8'h00;
im[4628]= 8'h03;
im[4629]= 8'h25;
im[4630]= 8'h84;
im[4631]= 8'hFA;
im[4632]= 8'h93;
im[4633]= 8'h15;
im[4634]= 8'h35;
im[4635]= 8'h00;
im[4636]= 8'h13;
im[4637]= 8'h05;
im[4638]= 8'h84;
im[4639]= 8'hFB;
im[4640]= 8'h33;
im[4641]= 8'h05;
im[4642]= 8'hB5;
im[4643]= 8'h00;
im[4644]= 8'h03;
im[4645]= 8'h26;
im[4646]= 8'h84;
im[4647]= 8'hF8;
im[4648]= 8'h83;
im[4649]= 8'h26;
im[4650]= 8'hC4;
im[4651]= 8'hF8;
im[4652]= 8'h6F;
im[4653]= 8'h00;
im[4654]= 8'h40;
im[4655]= 8'h00;
im[4656]= 8'h03;
im[4657]= 8'h25;
im[4658]= 8'h84;
im[4659]= 8'hFA;
im[4660]= 8'h13;
im[4661]= 8'h05;
im[4662]= 8'h15;
im[4663]= 8'h00;
im[4664]= 8'h23;
im[4665]= 8'h24;
im[4666]= 8'hA4;
im[4667]= 8'hFA;
im[4668]= 8'h6F;
im[4669]= 8'hF0;
im[4670]= 8'h9F;
im[4671]= 8'hFC;
im[4672]= 8'h23;
im[4673]= 8'h26;
im[4674]= 8'hA4;
im[4675]= 8'hFE;
im[4676]= 8'h23;
im[4677]= 8'h20;
im[4678]= 8'hA4;
im[4679]= 8'hF8;
im[4680]= 8'h23;
im[4681]= 8'h24;
im[4682]= 8'hA4;
im[4683]= 8'hFE;
im[4684]= 8'h23;
im[4685]= 8'h22;
im[4686]= 8'hB4;
im[4687]= 8'hFE;
im[4688]= 8'h23;
im[4689]= 8'h20;
im[4690]= 8'hA4;
im[4691]= 8'hFE;
im[4692]= 8'h23;
im[4693]= 8'h2E;
im[4694]= 8'hB4;
im[4695]= 8'hFC;
im[4696]= 8'h23;
im[4697]= 8'h2C;
im[4698]= 8'hA4;
im[4699]= 8'hFC;
im[4700]= 8'h23;
im[4701]= 8'h2A;
im[4702]= 8'hB4;
im[4703]= 8'hFC;
im[4704]= 8'h23;
im[4705]= 8'h28;
im[4706]= 8'hA4;
im[4707]= 8'hFC;
im[4708]= 8'h13;
im[4709]= 8'h05;
im[4710]= 8'hC4;
im[4711]= 8'hFA;
im[4712]= 8'h93;
im[4713]= 8'h05;
im[4714]= 8'h84;
im[4715]= 8'hFB;
im[4716]= 8'h03;
im[4717]= 8'h25;
im[4718]= 8'h04;
im[4719]= 8'hF8;
im[4720]= 8'h23;
im[4721]= 8'h24;
im[4722]= 8'hA4;
im[4723]= 8'hFA;
im[4724]= 8'h6F;
im[4725]= 8'h00;
im[4726]= 8'h40;
im[4727]= 8'h00;
im[4728]= 8'h03;
im[4729]= 8'h25;
im[4730]= 8'h84;
im[4731]= 8'hFA;
im[4732]= 8'h83;
im[4733]= 8'h25;
im[4734]= 8'hC4;
im[4735]= 8'hFA;
im[4736]= 8'h63;
im[4737]= 8'h5A;
im[4738]= 8'hB5;
im[4739]= 8'h02;
im[4740]= 8'h6F;
im[4741]= 8'h00;
im[4742]= 8'h40;
im[4743]= 8'h00;
im[4744]= 8'h03;
im[4745]= 8'h25;
im[4746]= 8'h84;
im[4747]= 8'hFA;
im[4748]= 8'h93;
im[4749]= 8'h15;
im[4750]= 8'h35;
im[4751]= 8'h00;
im[4752]= 8'h13;
im[4753]= 8'h05;
im[4754]= 8'h84;
im[4755]= 8'hFB;
im[4756]= 8'h33;
im[4757]= 8'h05;
im[4758]= 8'hB5;
im[4759]= 8'h00;
im[4760]= 8'h03;
im[4761]= 8'h26;
im[4762]= 8'h84;
im[4763]= 8'hF8;
im[4764]= 8'h83;
im[4765]= 8'h26;
im[4766]= 8'hC4;
im[4767]= 8'hF8;
im[4768]= 8'h6F;
im[4769]= 8'h00;
im[4770]= 8'h40;
im[4771]= 8'h00;
im[4772]= 8'h03;
im[4773]= 8'h25;
im[4774]= 8'h84;
im[4775]= 8'hFA;
im[4776]= 8'h13;
im[4777]= 8'h05;
im[4778]= 8'h15;
im[4779]= 8'h00;
im[4780]= 8'h23;
im[4781]= 8'h24;
im[4782]= 8'hA4;
im[4783]= 8'hFA;
im[4784]= 8'h6F;
im[4785]= 8'hF0;
im[4786]= 8'h9F;
im[4787]= 8'hFC;
im[4788]= 8'h23;
im[4789]= 8'h26;
im[4790]= 8'hA4;
im[4791]= 8'hFE;
im[4792]= 8'h23;
im[4793]= 8'h2E;
im[4794]= 8'hA4;
im[4795]= 8'hF6;
im[4796]= 8'h23;
im[4797]= 8'h24;
im[4798]= 8'hA4;
im[4799]= 8'hFE;
im[4800]= 8'h23;
im[4801]= 8'h22;
im[4802]= 8'hB4;
im[4803]= 8'hFE;
im[4804]= 8'h23;
im[4805]= 8'h20;
im[4806]= 8'hA4;
im[4807]= 8'hFE;
im[4808]= 8'h23;
im[4809]= 8'h2E;
im[4810]= 8'hB4;
im[4811]= 8'hFC;
im[4812]= 8'h23;
im[4813]= 8'h2C;
im[4814]= 8'hA4;
im[4815]= 8'hFC;
im[4816]= 8'h23;
im[4817]= 8'h2A;
im[4818]= 8'hB4;
im[4819]= 8'hFC;
im[4820]= 8'h23;
im[4821]= 8'h28;
im[4822]= 8'hA4;
im[4823]= 8'hFC;
im[4824]= 8'h13;
im[4825]= 8'h05;
im[4826]= 8'hC4;
im[4827]= 8'hFA;
im[4828]= 8'h93;
im[4829]= 8'h05;
im[4830]= 8'h84;
im[4831]= 8'hFB;
im[4832]= 8'h03;
im[4833]= 8'h25;
im[4834]= 8'hC4;
im[4835]= 8'hF7;
im[4836]= 8'h23;
im[4837]= 8'h24;
im[4838]= 8'hA4;
im[4839]= 8'hFA;
im[4840]= 8'h6F;
im[4841]= 8'h00;
im[4842]= 8'h40;
im[4843]= 8'h00;
im[4844]= 8'h03;
im[4845]= 8'h25;
im[4846]= 8'h84;
im[4847]= 8'hFA;
im[4848]= 8'h83;
im[4849]= 8'h25;
im[4850]= 8'hC4;
im[4851]= 8'hFA;
im[4852]= 8'h63;
im[4853]= 8'h5A;
im[4854]= 8'hB5;
im[4855]= 8'h02;
im[4856]= 8'h6F;
im[4857]= 8'h00;
im[4858]= 8'h40;
im[4859]= 8'h00;
im[4860]= 8'h03;
im[4861]= 8'h25;
im[4862]= 8'h84;
im[4863]= 8'hFA;
im[4864]= 8'h93;
im[4865]= 8'h15;
im[4866]= 8'h35;
im[4867]= 8'h00;
im[4868]= 8'h13;
im[4869]= 8'h05;
im[4870]= 8'h84;
im[4871]= 8'hFB;
im[4872]= 8'h33;
im[4873]= 8'h05;
im[4874]= 8'hB5;
im[4875]= 8'h00;
im[4876]= 8'h03;
im[4877]= 8'h26;
im[4878]= 8'h84;
im[4879]= 8'hF8;
im[4880]= 8'h83;
im[4881]= 8'h26;
im[4882]= 8'hC4;
im[4883]= 8'hF8;
im[4884]= 8'h6F;
im[4885]= 8'h00;
im[4886]= 8'h40;
im[4887]= 8'h00;
im[4888]= 8'h03;
im[4889]= 8'h25;
im[4890]= 8'h84;
im[4891]= 8'hFA;
im[4892]= 8'h13;
im[4893]= 8'h05;
im[4894]= 8'h15;
im[4895]= 8'h00;
im[4896]= 8'h23;
im[4897]= 8'h24;
im[4898]= 8'hA4;
im[4899]= 8'hFA;
im[4900]= 8'h6F;
im[4901]= 8'hF0;
im[4902]= 8'h9F;
im[4903]= 8'hFC;
im[4904]= 8'h23;
im[4905]= 8'h26;
im[4906]= 8'hB4;
im[4907]= 8'hFE;
im[4908]= 8'h23;
im[4909]= 8'h2C;
im[4910]= 8'hA4;
im[4911]= 8'hF6;
im[4912]= 8'h23;
im[4913]= 8'h24;
im[4914]= 8'hA4;
im[4915]= 8'hFE;
im[4916]= 8'h13;
im[4917]= 8'h06;
im[4918]= 8'h66;
im[4919]= 8'h66;
im[4920]= 8'h23;
im[4921]= 8'h22;
im[4922]= 8'hC4;
im[4923]= 8'hFE;
im[4924]= 8'h13;
im[4925]= 8'h06;
im[4926]= 8'h66;
im[4927]= 8'h66;
im[4928]= 8'h23;
im[4929]= 8'h20;
im[4930]= 8'hC4;
im[4931]= 8'hFE;
im[4932]= 8'h23;
im[4933]= 8'h2E;
im[4934]= 8'hB4;
im[4935]= 8'hFC;
im[4936]= 8'h23;
im[4937]= 8'h2C;
im[4938]= 8'hA4;
im[4939]= 8'hFC;
im[4940]= 8'h23;
im[4941]= 8'h2A;
im[4942]= 8'hB4;
im[4943]= 8'hFC;
im[4944]= 8'h23;
im[4945]= 8'h28;
im[4946]= 8'hA4;
im[4947]= 8'hFC;
im[4948]= 8'h13;
im[4949]= 8'h05;
im[4950]= 8'hC4;
im[4951]= 8'hFA;
im[4952]= 8'h93;
im[4953]= 8'h05;
im[4954]= 8'h84;
im[4955]= 8'hFB;
im[4956]= 8'h03;
im[4957]= 8'h25;
im[4958]= 8'h84;
im[4959]= 8'hF7;
im[4960]= 8'h23;
im[4961]= 8'h24;
im[4962]= 8'hA4;
im[4963]= 8'hFA;
im[4964]= 8'h6F;
im[4965]= 8'h00;
im[4966]= 8'h40;
im[4967]= 8'h00;
im[4968]= 8'h03;
im[4969]= 8'h25;
im[4970]= 8'h84;
im[4971]= 8'hFA;
im[4972]= 8'h83;
im[4973]= 8'h25;
im[4974]= 8'hC4;
im[4975]= 8'hFA;
im[4976]= 8'h63;
im[4977]= 8'h5A;
im[4978]= 8'hB5;
im[4979]= 8'h02;
im[4980]= 8'h6F;
im[4981]= 8'h00;
im[4982]= 8'h40;
im[4983]= 8'h00;
im[4984]= 8'h03;
im[4985]= 8'h25;
im[4986]= 8'h84;
im[4987]= 8'hFA;
im[4988]= 8'h93;
im[4989]= 8'h15;
im[4990]= 8'h35;
im[4991]= 8'h00;
im[4992]= 8'h13;
im[4993]= 8'h05;
im[4994]= 8'h84;
im[4995]= 8'hFB;
im[4996]= 8'h33;
im[4997]= 8'h05;
im[4998]= 8'hB5;
im[4999]= 8'h00;
im[5000]= 8'h03;
im[5001]= 8'h26;
im[5002]= 8'h84;
im[5003]= 8'hF8;
im[5004]= 8'h83;
im[5005]= 8'h26;
im[5006]= 8'hC4;
im[5007]= 8'hF8;
im[5008]= 8'h6F;
im[5009]= 8'h00;
im[5010]= 8'h40;
im[5011]= 8'h00;
im[5012]= 8'h03;
im[5013]= 8'h25;
im[5014]= 8'h84;
im[5015]= 8'hFA;
im[5016]= 8'h13;
im[5017]= 8'h05;
im[5018]= 8'h15;
im[5019]= 8'h00;
im[5020]= 8'h23;
im[5021]= 8'h24;
im[5022]= 8'hA4;
im[5023]= 8'hFA;
im[5024]= 8'h6F;
im[5025]= 8'hF0;
im[5026]= 8'h9F;
im[5027]= 8'hFC;
im[5028]= 8'h23;
im[5029]= 8'h26;
im[5030]= 8'hA4;
im[5031]= 8'hFE;
im[5032]= 8'h23;
im[5033]= 8'h2A;
im[5034]= 8'hA4;
im[5035]= 8'hF6;
im[5036]= 8'h23;
im[5037]= 8'h24;
im[5038]= 8'hA4;
im[5039]= 8'hFE;
im[5040]= 8'h93;
im[5041]= 8'h85;
im[5042]= 8'h45;
im[5043]= 8'hE1;
im[5044]= 8'h23;
im[5045]= 8'h22;
im[5046]= 8'hB4;
im[5047]= 8'hFE;
im[5048]= 8'h93;
im[5049]= 8'h85;
im[5050]= 8'hE5;
im[5051]= 8'h7A;
im[5052]= 8'h23;
im[5053]= 8'h20;
im[5054]= 8'hB4;
im[5055]= 8'hFE;
im[5056]= 8'h23;
im[5057]= 8'h2E;
im[5058]= 8'hB4;
im[5059]= 8'hFC;
im[5060]= 8'h23;
im[5061]= 8'h2C;
im[5062]= 8'hA4;
im[5063]= 8'hFC;
im[5064]= 8'h23;
im[5065]= 8'h2A;
im[5066]= 8'hB4;
im[5067]= 8'hFC;
im[5068]= 8'h23;
im[5069]= 8'h28;
im[5070]= 8'hA4;
im[5071]= 8'hFC;
im[5072]= 8'h13;
im[5073]= 8'h05;
im[5074]= 8'hC4;
im[5075]= 8'hFA;
im[5076]= 8'h93;
im[5077]= 8'h05;
im[5078]= 8'h84;
im[5079]= 8'hFB;
im[5080]= 8'h03;
im[5081]= 8'h25;
im[5082]= 8'h44;
im[5083]= 8'hF7;
im[5084]= 8'h23;
im[5085]= 8'h24;
im[5086]= 8'hA4;
im[5087]= 8'hFA;
im[5088]= 8'h6F;
im[5089]= 8'h00;
im[5090]= 8'h40;
im[5091]= 8'h00;
im[5092]= 8'h03;
im[5093]= 8'h25;
im[5094]= 8'h84;
im[5095]= 8'hFA;
im[5096]= 8'h83;
im[5097]= 8'h25;
im[5098]= 8'hC4;
im[5099]= 8'hFA;
im[5100]= 8'h63;
im[5101]= 8'h5A;
im[5102]= 8'hB5;
im[5103]= 8'h02;
im[5104]= 8'h6F;
im[5105]= 8'h00;
im[5106]= 8'h40;
im[5107]= 8'h00;
im[5108]= 8'h03;
im[5109]= 8'h25;
im[5110]= 8'h84;
im[5111]= 8'hFA;
im[5112]= 8'h93;
im[5113]= 8'h15;
im[5114]= 8'h35;
im[5115]= 8'h00;
im[5116]= 8'h13;
im[5117]= 8'h05;
im[5118]= 8'h84;
im[5119]= 8'hFB;
im[5120]= 8'h33;
im[5121]= 8'h05;
im[5122]= 8'hB5;
im[5123]= 8'h00;
im[5124]= 8'h03;
im[5125]= 8'h26;
im[5126]= 8'h84;
im[5127]= 8'hF8;
im[5128]= 8'h83;
im[5129]= 8'h26;
im[5130]= 8'hC4;
im[5131]= 8'hF8;
im[5132]= 8'h6F;
im[5133]= 8'h00;
im[5134]= 8'h40;
im[5135]= 8'h00;
im[5136]= 8'h03;
im[5137]= 8'h25;
im[5138]= 8'h84;
im[5139]= 8'hFA;
im[5140]= 8'h13;
im[5141]= 8'h05;
im[5142]= 8'h15;
im[5143]= 8'h00;
im[5144]= 8'h23;
im[5145]= 8'h24;
im[5146]= 8'hA4;
im[5147]= 8'hFA;
im[5148]= 8'h6F;
im[5149]= 8'hF0;
im[5150]= 8'h9F;
im[5151]= 8'hFC;
im[5152]= 8'h23;
im[5153]= 8'h26;
im[5154]= 8'hA4;
im[5155]= 8'hFE;
im[5156]= 8'h23;
im[5157]= 8'h28;
im[5158]= 8'hA4;
im[5159]= 8'hF6;
im[5160]= 8'h23;
im[5161]= 8'h24;
im[5162]= 8'hA4;
im[5163]= 8'hFE;
im[5164]= 8'h93;
im[5165]= 8'h85;
im[5166]= 8'h55;
im[5167]= 8'h8F;
im[5168]= 8'h23;
im[5169]= 8'h22;
im[5170]= 8'hB4;
im[5171]= 8'hFE;
im[5172]= 8'h93;
im[5173]= 8'h85;
im[5174]= 8'h95;
im[5175]= 8'hC2;
im[5176]= 8'h23;
im[5177]= 8'h20;
im[5178]= 8'hB4;
im[5179]= 8'hFE;
im[5180]= 8'h23;
im[5181]= 8'h2E;
im[5182]= 8'hB4;
im[5183]= 8'hFC;
im[5184]= 8'h23;
im[5185]= 8'h2C;
im[5186]= 8'hA4;
im[5187]= 8'hFC;
im[5188]= 8'h13;
im[5189]= 8'h05;
im[5190]= 8'h95;
im[5191]= 8'h99;
im[5192]= 8'h23;
im[5193]= 8'h2A;
im[5194]= 8'hA4;
im[5195]= 8'hFC;
im[5196]= 8'h13;
im[5197]= 8'h05;
im[5198]= 8'hA5;
im[5199]= 8'h99;
im[5200]= 8'h23;
im[5201]= 8'h28;
im[5202]= 8'hA4;
im[5203]= 8'hFC;
im[5204]= 8'h13;
im[5205]= 8'h05;
im[5206]= 8'hC4;
im[5207]= 8'hFA;
im[5208]= 8'h93;
im[5209]= 8'h05;
im[5210]= 8'h84;
im[5211]= 8'hFB;
im[5212]= 8'h03;
im[5213]= 8'h25;
im[5214]= 8'h04;
im[5215]= 8'hF7;
im[5216]= 8'h23;
im[5217]= 8'h24;
im[5218]= 8'hA4;
im[5219]= 8'hFA;
im[5220]= 8'h6F;
im[5221]= 8'h00;
im[5222]= 8'h40;
im[5223]= 8'h00;
im[5224]= 8'h03;
im[5225]= 8'h25;
im[5226]= 8'h84;
im[5227]= 8'hFA;
im[5228]= 8'h83;
im[5229]= 8'h25;
im[5230]= 8'hC4;
im[5231]= 8'hFA;
im[5232]= 8'h63;
im[5233]= 8'h5A;
im[5234]= 8'hB5;
im[5235]= 8'h02;
im[5236]= 8'h6F;
im[5237]= 8'h00;
im[5238]= 8'h40;
im[5239]= 8'h00;
im[5240]= 8'h03;
im[5241]= 8'h25;
im[5242]= 8'h84;
im[5243]= 8'hFA;
im[5244]= 8'h93;
im[5245]= 8'h15;
im[5246]= 8'h35;
im[5247]= 8'h00;
im[5248]= 8'h13;
im[5249]= 8'h05;
im[5250]= 8'h84;
im[5251]= 8'hFB;
im[5252]= 8'h33;
im[5253]= 8'h05;
im[5254]= 8'hB5;
im[5255]= 8'h00;
im[5256]= 8'h03;
im[5257]= 8'h26;
im[5258]= 8'h84;
im[5259]= 8'hF8;
im[5260]= 8'h83;
im[5261]= 8'h26;
im[5262]= 8'hC4;
im[5263]= 8'hF8;
im[5264]= 8'h6F;
im[5265]= 8'h00;
im[5266]= 8'h40;
im[5267]= 8'h00;
im[5268]= 8'h03;
im[5269]= 8'h25;
im[5270]= 8'h84;
im[5271]= 8'hFA;
im[5272]= 8'h13;
im[5273]= 8'h05;
im[5274]= 8'h15;
im[5275]= 8'h00;
im[5276]= 8'h23;
im[5277]= 8'h24;
im[5278]= 8'hA4;
im[5279]= 8'hFA;
im[5280]= 8'h6F;
im[5281]= 8'hF0;
im[5282]= 8'h9F;
im[5283]= 8'hFC;
im[5284]= 8'h23;
im[5285]= 8'h26;
im[5286]= 8'hA4;
im[5287]= 8'hFE;
im[5288]= 8'h23;
im[5289]= 8'h26;
im[5290]= 8'hA4;
im[5291]= 8'hF6;
im[5292]= 8'h23;
im[5293]= 8'h24;
im[5294]= 8'hA4;
im[5295]= 8'hFE;
im[5296]= 8'h93;
im[5297]= 8'h85;
im[5298]= 8'hA5;
im[5299]= 8'h70;
im[5300]= 8'h23;
im[5301]= 8'h22;
im[5302]= 8'hB4;
im[5303]= 8'hFE;
im[5304]= 8'h93;
im[5305]= 8'h85;
im[5306]= 8'h75;
im[5307]= 8'h3D;
im[5308]= 8'h23;
im[5309]= 8'h20;
im[5310]= 8'hB4;
im[5311]= 8'hFE;
im[5312]= 8'h23;
im[5313]= 8'h2E;
im[5314]= 8'hB4;
im[5315]= 8'hFC;
im[5316]= 8'h23;
im[5317]= 8'h2C;
im[5318]= 8'hA4;
im[5319]= 8'hFC;
im[5320]= 8'h23;
im[5321]= 8'h2A;
im[5322]= 8'hB4;
im[5323]= 8'hFC;
im[5324]= 8'h23;
im[5325]= 8'h28;
im[5326]= 8'hA4;
im[5327]= 8'hFC;
im[5328]= 8'h13;
im[5329]= 8'h05;
im[5330]= 8'hC4;
im[5331]= 8'hFA;
im[5332]= 8'h93;
im[5333]= 8'h05;
im[5334]= 8'h84;
im[5335]= 8'hFB;
im[5336]= 8'h03;
im[5337]= 8'h25;
im[5338]= 8'hC4;
im[5339]= 8'hF6;
im[5340]= 8'h23;
im[5341]= 8'h24;
im[5342]= 8'hA4;
im[5343]= 8'hFA;
im[5344]= 8'h6F;
im[5345]= 8'h00;
im[5346]= 8'h40;
im[5347]= 8'h00;
im[5348]= 8'h03;
im[5349]= 8'h25;
im[5350]= 8'h84;
im[5351]= 8'hFA;
im[5352]= 8'h83;
im[5353]= 8'h25;
im[5354]= 8'hC4;
im[5355]= 8'hFA;
im[5356]= 8'h63;
im[5357]= 8'h5A;
im[5358]= 8'hB5;
im[5359]= 8'h02;
im[5360]= 8'h6F;
im[5361]= 8'h00;
im[5362]= 8'h40;
im[5363]= 8'h00;
im[5364]= 8'h03;
im[5365]= 8'h25;
im[5366]= 8'h84;
im[5367]= 8'hFA;
im[5368]= 8'h93;
im[5369]= 8'h15;
im[5370]= 8'h35;
im[5371]= 8'h00;
im[5372]= 8'h13;
im[5373]= 8'h05;
im[5374]= 8'h84;
im[5375]= 8'hFB;
im[5376]= 8'h33;
im[5377]= 8'h05;
im[5378]= 8'hB5;
im[5379]= 8'h00;
im[5380]= 8'h03;
im[5381]= 8'h26;
im[5382]= 8'h84;
im[5383]= 8'hF8;
im[5384]= 8'h83;
im[5385]= 8'h26;
im[5386]= 8'hC4;
im[5387]= 8'hF8;
im[5388]= 8'h6F;
im[5389]= 8'h00;
im[5390]= 8'h40;
im[5391]= 8'h00;
im[5392]= 8'h03;
im[5393]= 8'h25;
im[5394]= 8'h84;
im[5395]= 8'hFA;
im[5396]= 8'h13;
im[5397]= 8'h05;
im[5398]= 8'h15;
im[5399]= 8'h00;
im[5400]= 8'h23;
im[5401]= 8'h24;
im[5402]= 8'hA4;
im[5403]= 8'hFA;
im[5404]= 8'h6F;
im[5405]= 8'hF0;
im[5406]= 8'h9F;
im[5407]= 8'hFC;
im[5408]= 8'h23;
im[5409]= 8'h26;
im[5410]= 8'hA4;
im[5411]= 8'hFE;
im[5412]= 8'h23;
im[5413]= 8'h24;
im[5414]= 8'hA4;
im[5415]= 8'hF6;
im[5416]= 8'h23;
im[5417]= 8'h24;
im[5418]= 8'hA4;
im[5419]= 8'hFE;
im[5420]= 8'h93;
im[5421]= 8'h85;
im[5422]= 8'h35;
im[5423]= 8'h33;
im[5424]= 8'h23;
im[5425]= 8'h22;
im[5426]= 8'hB4;
im[5427]= 8'hFE;
im[5428]= 8'h93;
im[5429]= 8'h85;
im[5430]= 8'h35;
im[5431]= 8'h33;
im[5432]= 8'h23;
im[5433]= 8'h20;
im[5434]= 8'hB4;
im[5435]= 8'hFE;
im[5436]= 8'h13;
im[5437]= 8'h06;
im[5438]= 8'h36;
im[5439]= 8'h33;
im[5440]= 8'h23;
im[5441]= 8'h2E;
im[5442]= 8'hC4;
im[5443]= 8'hFC;
im[5444]= 8'h23;
im[5445]= 8'h2C;
im[5446]= 8'hB4;
im[5447]= 8'hFC;
im[5448]= 8'h23;
im[5449]= 8'h2A;
im[5450]= 8'hB4;
im[5451]= 8'hFC;
im[5452]= 8'h23;
im[5453]= 8'h28;
im[5454]= 8'hA4;
im[5455]= 8'hFC;
im[5456]= 8'h13;
im[5457]= 8'h05;
im[5458]= 8'hC4;
im[5459]= 8'hFA;
im[5460]= 8'h93;
im[5461]= 8'h05;
im[5462]= 8'h84;
im[5463]= 8'hFB;
im[5464]= 8'h03;
im[5465]= 8'h25;
im[5466]= 8'h84;
im[5467]= 8'hF6;
im[5468]= 8'h23;
im[5469]= 8'h24;
im[5470]= 8'hA4;
im[5471]= 8'hFA;
im[5472]= 8'h6F;
im[5473]= 8'h00;
im[5474]= 8'h40;
im[5475]= 8'h00;
im[5476]= 8'h03;
im[5477]= 8'h25;
im[5478]= 8'h84;
im[5479]= 8'hFA;
im[5480]= 8'h83;
im[5481]= 8'h25;
im[5482]= 8'hC4;
im[5483]= 8'hFA;
im[5484]= 8'h63;
im[5485]= 8'h5A;
im[5486]= 8'hB5;
im[5487]= 8'h02;
im[5488]= 8'h6F;
im[5489]= 8'h00;
im[5490]= 8'h40;
im[5491]= 8'h00;
im[5492]= 8'h03;
im[5493]= 8'h25;
im[5494]= 8'h84;
im[5495]= 8'hFA;
im[5496]= 8'h93;
im[5497]= 8'h15;
im[5498]= 8'h35;
im[5499]= 8'h00;
im[5500]= 8'h13;
im[5501]= 8'h05;
im[5502]= 8'h84;
im[5503]= 8'hFB;
im[5504]= 8'h33;
im[5505]= 8'h05;
im[5506]= 8'hB5;
im[5507]= 8'h00;
im[5508]= 8'h03;
im[5509]= 8'h26;
im[5510]= 8'h84;
im[5511]= 8'hF8;
im[5512]= 8'h83;
im[5513]= 8'h26;
im[5514]= 8'hC4;
im[5515]= 8'hF8;
im[5516]= 8'h6F;
im[5517]= 8'h00;
im[5518]= 8'h40;
im[5519]= 8'h00;
im[5520]= 8'h03;
im[5521]= 8'h25;
im[5522]= 8'h84;
im[5523]= 8'hFA;
im[5524]= 8'h13;
im[5525]= 8'h05;
im[5526]= 8'h15;
im[5527]= 8'h00;
im[5528]= 8'h23;
im[5529]= 8'h24;
im[5530]= 8'hA4;
im[5531]= 8'hFA;
im[5532]= 8'h6F;
im[5533]= 8'hF0;
im[5534]= 8'h9F;
im[5535]= 8'hFC;
im[5536]= 8'h23;
im[5537]= 8'h26;
im[5538]= 8'hA4;
im[5539]= 8'hFE;
im[5540]= 8'h23;
im[5541]= 8'h24;
im[5542]= 8'hA4;
im[5543]= 8'hFE;
im[5544]= 8'h6F;
im[5545]= 8'h00;
im[5546]= 8'h40;
im[5547]= 8'h00;
im[5548]= 8'h6F;
im[5549]= 8'h00;
im[5550]= 8'h40;
im[5551]= 8'h00;
im[5552]= 8'h23;
im[5553]= 8'h22;
im[5554]= 8'hA4;
im[5555]= 8'hFE;
im[5556]= 8'h23;
im[5557]= 8'h20;
im[5558]= 8'hA4;
im[5559]= 8'hFE;
im[5560]= 8'h6F;
im[5561]= 8'h00;
im[5562]= 8'h40;
im[5563]= 8'h00;
im[5564]= 8'h6F;
im[5565]= 8'h00;
im[5566]= 8'h40;
im[5567]= 8'h00;
im[5568]= 8'h23;
im[5569]= 8'h2E;
im[5570]= 8'hA4;
im[5571]= 8'hFC;
im[5572]= 8'h23;
im[5573]= 8'h2C;
im[5574]= 8'hA4;
im[5575]= 8'hFC;
im[5576]= 8'h6F;
im[5577]= 8'h00;
im[5578]= 8'h40;
im[5579]= 8'h00;
im[5580]= 8'h6F;
im[5581]= 8'h00;
im[5582]= 8'h40;
im[5583]= 8'h00;
im[5584]= 8'h23;
im[5585]= 8'h2A;
im[5586]= 8'hA4;
im[5587]= 8'hFC;
im[5588]= 8'h23;
im[5589]= 8'h28;
im[5590]= 8'hA4;
im[5591]= 8'hFC;
im[5592]= 8'h6F;
im[5593]= 8'h00;
im[5594]= 8'h40;
im[5595]= 8'h00;
im[5596]= 8'h6F;
im[5597]= 8'h00;
im[5598]= 8'h40;
im[5599]= 8'h00;
im[5600]= 8'h13;
im[5601]= 8'h05;
im[5602]= 8'hC4;
im[5603]= 8'hFA;
im[5604]= 8'h93;
im[5605]= 8'h05;
im[5606]= 8'h84;
im[5607]= 8'hFB;
im[5608]= 8'h23;
im[5609]= 8'h24;
im[5610]= 8'hA4;
im[5611]= 8'hFA;
im[5612]= 8'h6F;
im[5613]= 8'h00;
im[5614]= 8'h40;
im[5615]= 8'h00;
im[5616]= 8'h03;
im[5617]= 8'h25;
im[5618]= 8'h84;
im[5619]= 8'hFA;
im[5620]= 8'h83;
im[5621]= 8'h25;
im[5622]= 8'hC4;
im[5623]= 8'hFA;
im[5624]= 8'h63;
im[5625]= 8'h5A;
im[5626]= 8'hB5;
im[5627]= 8'h02;
im[5628]= 8'h6F;
im[5629]= 8'h00;
im[5630]= 8'h40;
im[5631]= 8'h00;
im[5632]= 8'h03;
im[5633]= 8'h25;
im[5634]= 8'h84;
im[5635]= 8'hFA;
im[5636]= 8'h93;
im[5637]= 8'h15;
im[5638]= 8'h35;
im[5639]= 8'h00;
im[5640]= 8'h13;
im[5641]= 8'h05;
im[5642]= 8'h84;
im[5643]= 8'hFB;
im[5644]= 8'h33;
im[5645]= 8'h05;
im[5646]= 8'hB5;
im[5647]= 8'h00;
im[5648]= 8'h03;
im[5649]= 8'h26;
im[5650]= 8'h84;
im[5651]= 8'hF8;
im[5652]= 8'h83;
im[5653]= 8'h26;
im[5654]= 8'hC4;
im[5655]= 8'hF8;
im[5656]= 8'h6F;
im[5657]= 8'h00;
im[5658]= 8'h40;
im[5659]= 8'h00;
im[5660]= 8'h03;
im[5661]= 8'h25;
im[5662]= 8'h84;
im[5663]= 8'hFA;
im[5664]= 8'h13;
im[5665]= 8'h05;
im[5666]= 8'h15;
im[5667]= 8'h00;
im[5668]= 8'h23;
im[5669]= 8'h24;
im[5670]= 8'hA4;
im[5671]= 8'hFA;
im[5672]= 8'h6F;
im[5673]= 8'hF0;
im[5674]= 8'h9F;
im[5675]= 8'hFC;
im[5676]= 8'h6F;
im[5677]= 8'h00;
im[5678]= 8'h40;
im[5679]= 8'h00;
im[5680]= 8'h6F;
im[5681]= 8'hF0;
im[5682]= 8'hDF;
im[5683]= 8'hFA;
im[5684]= 8'h6F;
im[5685]= 8'h00;
im[5686]= 8'h40;
im[5687]= 8'h00;
im[5688]= 8'h6F;
im[5689]= 8'hF0;
im[5690]= 8'h5F;
im[5691]= 8'hF9;
im[5692]= 8'h6F;
im[5693]= 8'h00;
im[5694]= 8'h40;
im[5695]= 8'h00;
im[5696]= 8'h6F;
im[5697]= 8'hF0;
im[5698]= 8'hDF;
im[5699]= 8'hF7;
im[5700]= 8'h6F;
im[5701]= 8'h00;
im[5702]= 8'h40;
im[5703]= 8'h00;
im[5704]= 8'h6F;
im[5705]= 8'hF0;
im[5706]= 8'h5F;
im[5707]= 8'hF6;
im[5708]= 8'h23;
im[5709]= 8'h24;
im[5710]= 8'hA4;
im[5711]= 8'hFA;
im[5712]= 8'h6F;
im[5713]= 8'h00;
im[5714]= 8'h40;
im[5715]= 8'h00;
im[5716]= 8'h83;
im[5717]= 8'h25;
im[5718]= 8'h84;
im[5719]= 8'hFA;
im[5720]= 8'h13;
im[5721]= 8'h05;
im[5722]= 8'hF5;
im[5723]= 8'h69;
im[5724]= 8'h63;
im[5725]= 8'h46;
im[5726]= 8'hB5;
im[5727]= 8'h02;
im[5728]= 8'h6F;
im[5729]= 8'h00;
im[5730]= 8'h40;
im[5731]= 8'h00;
im[5732]= 8'h03;
im[5733]= 8'h25;
im[5734]= 8'h84;
im[5735]= 8'hFA;
im[5736]= 8'h93;
im[5737]= 8'h05;
im[5738]= 8'h84;
im[5739]= 8'hF9;
im[5740]= 8'h83;
im[5741]= 8'h25;
im[5742]= 8'h84;
im[5743]= 8'hFA;
im[5744]= 8'h03;
im[5745]= 8'h26;
im[5746]= 8'h84;
im[5747]= 8'hF9;
im[5748]= 8'h6F;
im[5749]= 8'h00;
im[5750]= 8'h40;
im[5751]= 8'h00;
im[5752]= 8'h03;
im[5753]= 8'h25;
im[5754]= 8'h84;
im[5755]= 8'hFA;
im[5756]= 8'h13;
im[5757]= 8'h05;
im[5758]= 8'h25;
im[5759]= 8'h00;
im[5760]= 8'h23;
im[5761]= 8'h24;
im[5762]= 8'hA4;
im[5763]= 8'hFA;
im[5764]= 8'h6F;
im[5765]= 8'hF0;
im[5766]= 8'h1F;
im[5767]= 8'hFD;
im[5768]= 8'h13;
im[5769]= 8'h05;
im[5770]= 8'h95;
im[5771]= 8'h16;
im[5772]= 8'h23;
im[5773]= 8'h22;
im[5774]= 8'hA4;
im[5775]= 8'hFA;
im[5776]= 8'h6F;
im[5777]= 8'h00;
im[5778]= 8'h40;
im[5779]= 8'h00;
im[5780]= 8'h83;
im[5781]= 8'h25;
im[5782]= 8'h44;
im[5783]= 8'hFA;
im[5784]= 8'h13;
im[5785]= 8'h05;
im[5786]= 8'h85;
im[5787]= 8'h16;
im[5788]= 8'h63;
im[5789]= 8'h66;
im[5790]= 8'hB5;
im[5791]= 8'h02;
im[5792]= 8'h6F;
im[5793]= 8'h00;
im[5794]= 8'h40;
im[5795]= 8'h00;
im[5796]= 8'h03;
im[5797]= 8'h25;
im[5798]= 8'h44;
im[5799]= 8'hFA;
im[5800]= 8'h93;
im[5801]= 8'h05;
im[5802]= 8'h84;
im[5803]= 8'hF9;
im[5804]= 8'h83;
im[5805]= 8'h25;
im[5806]= 8'h44;
im[5807]= 8'hFA;
im[5808]= 8'h03;
im[5809]= 8'h26;
im[5810]= 8'h84;
im[5811]= 8'hF9;
im[5812]= 8'h6F;
im[5813]= 8'h00;
im[5814]= 8'h40;
im[5815]= 8'h00;
im[5816]= 8'h03;
im[5817]= 8'h25;
im[5818]= 8'h44;
im[5819]= 8'hFA;
im[5820]= 8'h13;
im[5821]= 8'h05;
im[5822]= 8'h15;
im[5823]= 8'h00;
im[5824]= 8'h23;
im[5825]= 8'h22;
im[5826]= 8'hA4;
im[5827]= 8'hFA;
im[5828]= 8'h6F;
im[5829]= 8'hF0;
im[5830]= 8'h1F;
im[5831]= 8'hFD;
im[5832]= 8'h23;
im[5833]= 8'h2A;
im[5834]= 8'hA4;
im[5835]= 8'hFA;
im[5836]= 8'h23;
im[5837]= 8'h28;
im[5838]= 8'hA4;
im[5839]= 8'hFA;
im[5840]= 8'h6F;
im[5841]= 8'h00;
im[5842]= 8'h40;
im[5843]= 8'h00;
im[5844]= 8'h6F;
im[5845]= 8'h00;
im[5846]= 8'h40;
im[5847]= 8'h00;
im[5848]= 8'h03;
im[5849]= 8'h27;
im[5850]= 8'h84;
im[5851]= 8'hF8;
im[5852]= 8'h83;
im[5853]= 8'h27;
im[5854]= 8'hC4;
im[5855]= 8'hF8;
im[5856]= 8'h03;
im[5857]= 8'h26;
im[5858]= 8'h84;
im[5859]= 8'hF8;
im[5860]= 8'h83;
im[5861]= 8'h26;
im[5862]= 8'hC4;
im[5863]= 8'hF8;
im[5864]= 8'h6F;
im[5865]= 8'h00;
im[5866]= 8'h40;
im[5867]= 8'h00;
im[5868]= 8'h6F;
im[5869]= 8'hF0;
im[5870]= 8'h9F;
im[5871]= 8'hFE;
im[5872]= 8'h23;
im[5873]= 8'h2A;
im[5874]= 8'hA4;
im[5875]= 8'hFA;
im[5876]= 8'h23;
im[5877]= 8'h28;
im[5878]= 8'hA4;
im[5879]= 8'hFA;
im[5880]= 8'h6F;
im[5881]= 8'h00;
im[5882]= 8'h40;
im[5883]= 8'h00;
im[5884]= 8'h6F;
im[5885]= 8'h00;
im[5886]= 8'h40;
im[5887]= 8'h00;
im[5888]= 8'h03;
im[5889]= 8'h27;
im[5890]= 8'h84;
im[5891]= 8'hF8;
im[5892]= 8'h83;
im[5893]= 8'h27;
im[5894]= 8'hC4;
im[5895]= 8'hF8;
im[5896]= 8'h03;
im[5897]= 8'h26;
im[5898]= 8'h84;
im[5899]= 8'hF8;
im[5900]= 8'h83;
im[5901]= 8'h26;
im[5902]= 8'hC4;
im[5903]= 8'hF8;
im[5904]= 8'h6F;
im[5905]= 8'h00;
im[5906]= 8'h40;
im[5907]= 8'h00;
im[5908]= 8'h6F;
im[5909]= 8'hF0;
im[5910]= 8'h9F;
im[5911]= 8'hFE;
im[5912]= 8'h03;
im[5913]= 8'h24;
im[5914]= 8'h81;
im[5915]= 8'h0B;
im[5916]= 8'h83;
im[5917]= 8'h20;
im[5918]= 8'hC1;
im[5919]= 8'h0B;
im[5920]= 8'h13;
im[5921]= 8'h01;
im[5922]= 8'h01;
im[5923]= 8'h0C;

end
always @ (*) begin //reSading pc to output instruction
data_out={im[PCn+3],im[PCn+2],im[PCn+1],im[PCn]};
//data_out=#5 {im[PCn+3],im[PCn+2],im[PCn+1],im[PCn]};
end

endmodule 

module add4(PC,PC4); //incrementing PC by 4
//input clk;
parameter PCSIZE=16;

input [PCSIZE-1:0] PC;
output  [PCSIZE-1:0] PC4;

assign PC4=PC+16'd4;

endmodule 